module mult_32b_5s ( 
input [32-1:0] a,
input [32-1:0] b,
output [2*32-1:0] r
);

// Target value:1157
wire [59:0] P;
wire [59:0] G;

// 4 normal LUT
LUT6_2 #(
.INIT(64'h78887888C0C0C0C0)
) LUT6_2_inst_f0 (
.O6(r[1]),
.O5(r[0]),
.I0(b[1]),
.I1(a[0]),
.I2(b[0]),
.I3(a[1]),
.I4(1'b1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h47777888B8887888)
) LUT6_2_inst_f1 (
.O6(r[2]),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

LUT6_2 #(
.INIT(64'hF8888000C0008000)
) LUT6_2_inst_f2 (
.O6(C1),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

LUT6_2 #(
.INIT(64'h8000000000000000)
) LUT6_2_inst_f3 (
.O6(C0),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

/////////STEP0----ORDER0////////////

wire p_s0_o0_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o0_t0_z0_v0 (
.O6(p_s0_o0_0),
.O5(),
.I0(a[3]),
.I1(b[0]),
.I2(a[2]),
.I3(b[1]),
.I4(a[1]),
.I5(b[2]));

wire p_s0_o1_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o0_t0_z1_v0 (
.O6(p_s0_o1_0),
.O5(),
.I0(a[3]),
.I1(b[0]),
.I2(a[2]),
.I3(b[1]),
.I4(a[1]),
.I5(b[2]));

/////////STEP0----ORDER1////////////

/////////STEP0----ORDER2////////////

/////////STEP0----ORDER3////////////

wire p_s0_o3_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o3_t1_z0_v0 (
.O6(p_s0_o3_0),
.O5(),
.I0(a[6]),
.I1(b[0]),
.I2(a[5]),
.I3(b[1]),
.I4(a[4]),
.I5(b[2]));

wire p_s0_o4_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o3_t1_z1_v0 (
.O6(p_s0_o4_0),
.O5(),
.I0(a[6]),
.I1(b[0]),
.I2(a[5]),
.I3(b[1]),
.I4(a[4]),
.I5(b[2]));

/////////STEP0----ORDER4////////////

wire p_s0_o4_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o4_t2_z0_v0 (
.O6(p_s0_o4_1),
.O5(),
.I0(a[7]),
.I1(b[0]),
.I2(a[6]),
.I3(b[1]),
.I4(a[5]),
.I5(b[2]));

wire p_s0_o5_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o4_t2_z1_v0 (
.O6(p_s0_o5_0),
.O5(),
.I0(a[7]),
.I1(b[0]),
.I2(a[6]),
.I3(b[1]),
.I4(a[5]),
.I5(b[2]));

/////////STEP0----ORDER5////////////

/////////STEP0----ORDER6////////////

/////////STEP0----ORDER7////////////

wire p_s0_o7_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o7_t3_z0_v0 (
.O6(p_s0_o7_0),
.O5(),
.I0(a[10]),
.I1(b[0]),
.I2(a[9]),
.I3(b[1]),
.I4(a[8]),
.I5(b[2]));

wire p_s0_o8_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o7_t3_z1_v0 (
.O6(p_s0_o8_0),
.O5(),
.I0(a[10]),
.I1(b[0]),
.I2(a[9]),
.I3(b[1]),
.I4(a[8]),
.I5(b[2]));

wire p_s0_o7_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o7_t3_z0_v1 (
.O6(p_s0_o7_1),
.O5(),
.I0(a[7]),
.I1(b[3]),
.I2(a[6]),
.I3(b[4]),
.I4(a[5]),
.I5(b[5]));

wire p_s0_o8_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o7_t3_z1_v1 (
.O6(p_s0_o8_1),
.O5(),
.I0(a[7]),
.I1(b[3]),
.I2(a[6]),
.I3(b[4]),
.I4(a[5]),
.I5(b[5]));

/////////STEP0----ORDER8////////////

/////////STEP0----ORDER9////////////

wire p_s0_o9_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o9_t4_z0_v0 (
.O6(p_s0_o9_0),
.O5(),
.I0(a[12]),
.I1(b[0]),
.I2(a[11]),
.I3(b[1]),
.I4(a[10]),
.I5(b[2]));

wire p_s0_o10_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o9_t4_z1_v0 (
.O6(p_s0_o10_0),
.O5(),
.I0(a[12]),
.I1(b[0]),
.I2(a[11]),
.I3(b[1]),
.I4(a[10]),
.I5(b[2]));

/////////STEP0----ORDER10////////////

wire p_s0_o10_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o10_t5_z0_v0 (
.O6(p_s0_o10_1),
.O5(),
.I0(a[13]),
.I1(b[0]),
.I2(a[12]),
.I3(b[1]),
.I4(a[11]),
.I5(b[2]));

wire p_s0_o11_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o10_t5_z1_v0 (
.O6(p_s0_o11_0),
.O5(),
.I0(a[13]),
.I1(b[0]),
.I2(a[12]),
.I3(b[1]),
.I4(a[11]),
.I5(b[2]));

wire p_s0_o10_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o10_t5_z0_v1 (
.O6(p_s0_o10_2),
.O5(),
.I0(a[10]),
.I1(b[3]),
.I2(a[9]),
.I3(b[4]),
.I4(a[8]),
.I5(b[5]));

wire p_s0_o11_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o10_t5_z1_v1 (
.O6(p_s0_o11_1),
.O5(),
.I0(a[10]),
.I1(b[3]),
.I2(a[9]),
.I3(b[4]),
.I4(a[8]),
.I5(b[5]));

/////////STEP0----ORDER11////////////

wire p_s0_o11_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o11_t6_z0_v0 (
.O6(p_s0_o11_2),
.O5(),
.I0(a[14]),
.I1(b[0]),
.I2(a[13]),
.I3(b[1]),
.I4(a[12]),
.I5(b[2]));

wire p_s0_o12_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o11_t6_z1_v0 (
.O6(p_s0_o12_0),
.O5(),
.I0(a[14]),
.I1(b[0]),
.I2(a[13]),
.I3(b[1]),
.I4(a[12]),
.I5(b[2]));

wire p_s0_o12_1;
wire p_s0_o11_3;
LUT6_2 #(
.INIT(64'h8000800078887888)
) LUT6_2_inst_s0_o11_t46_z0_v0 (
.O6(p_s0_o12_1),
.O5(p_s0_o11_3),
.I0(a[11]),
.I1(b[3]),
.I2(a[10]),
.I3(b[4]),
.I4(1'b0),
.I5(1'b1));

/////////STEP0----ORDER12////////////

wire p_s0_o13_0;
wire p_s0_o12_2;
LUT6_2 #(
.INIT(64'h8000800078887888)
) LUT6_2_inst_s0_o12_t47_z0_v0 (
.O6(p_s0_o13_0),
.O5(p_s0_o12_2),
.I0(a[15]),
.I1(b[0]),
.I2(a[14]),
.I3(b[1]),
.I4(1'b0),
.I5(1'b1));

/////////STEP0----ORDER13////////////

wire p_s0_o13_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o13_t7_z0_v0 (
.O6(p_s0_o13_1),
.O5(),
.I0(a[16]),
.I1(b[0]),
.I2(a[15]),
.I3(b[1]),
.I4(a[14]),
.I5(b[2]));

wire p_s0_o14_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o13_t7_z1_v0 (
.O6(p_s0_o14_0),
.O5(),
.I0(a[16]),
.I1(b[0]),
.I2(a[15]),
.I3(b[1]),
.I4(a[14]),
.I5(b[2]));

wire p_s0_o13_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o13_t7_z0_v1 (
.O6(p_s0_o13_2),
.O5(),
.I0(a[13]),
.I1(b[3]),
.I2(a[12]),
.I3(b[4]),
.I4(a[11]),
.I5(b[5]));

wire p_s0_o14_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o13_t7_z1_v1 (
.O6(p_s0_o14_1),
.O5(),
.I0(a[13]),
.I1(b[3]),
.I2(a[12]),
.I3(b[4]),
.I4(a[11]),
.I5(b[5]));

wire p_s0_o13_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o13_t7_z0_v2 (
.O6(p_s0_o13_3),
.O5(),
.I0(a[10]),
.I1(b[6]),
.I2(a[9]),
.I3(b[7]),
.I4(a[8]),
.I5(b[8]));

wire p_s0_o14_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o13_t7_z1_v2 (
.O6(p_s0_o14_2),
.O5(),
.I0(a[10]),
.I1(b[6]),
.I2(a[9]),
.I3(b[7]),
.I4(a[8]),
.I5(b[8]));

wire p_s0_o13_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o13_t7_z0_v3 (
.O6(p_s0_o13_4),
.O5(),
.I0(a[7]),
.I1(b[9]),
.I2(a[6]),
.I3(b[10]),
.I4(a[5]),
.I5(b[11]));

wire p_s0_o14_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o13_t7_z1_v3 (
.O6(p_s0_o14_3),
.O5(),
.I0(a[7]),
.I1(b[9]),
.I2(a[6]),
.I3(b[10]),
.I4(a[5]),
.I5(b[11]));

wire p_s0_o13_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o13_t7_z0_v4 (
.O6(p_s0_o13_5),
.O5(),
.I0(a[4]),
.I1(b[12]),
.I2(a[3]),
.I3(b[13]),
.I4(a[2]),
.I5(b[14]));

wire p_s0_o14_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o13_t7_z1_v4 (
.O6(p_s0_o14_4),
.O5(),
.I0(a[4]),
.I1(b[12]),
.I2(a[3]),
.I3(b[13]),
.I4(a[2]),
.I5(b[14]));

/////////STEP0----ORDER14////////////

wire p_s0_o14_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o14_t8_z0_v0 (
.O6(p_s0_o14_5),
.O5(),
.I0(a[17]),
.I1(b[0]),
.I2(a[16]),
.I3(b[1]),
.I4(a[15]),
.I5(b[2]));

wire p_s0_o15_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o14_t8_z1_v0 (
.O6(p_s0_o15_0),
.O5(),
.I0(a[17]),
.I1(b[0]),
.I2(a[16]),
.I3(b[1]),
.I4(a[15]),
.I5(b[2]));

wire p_s0_o14_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o14_t8_z0_v1 (
.O6(p_s0_o14_6),
.O5(),
.I0(a[14]),
.I1(b[3]),
.I2(a[13]),
.I3(b[4]),
.I4(a[12]),
.I5(b[5]));

wire p_s0_o15_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o14_t8_z1_v1 (
.O6(p_s0_o15_1),
.O5(),
.I0(a[14]),
.I1(b[3]),
.I2(a[13]),
.I3(b[4]),
.I4(a[12]),
.I5(b[5]));

/////////STEP0----ORDER15////////////

wire p_s0_o15_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o15_t9_z0_v0 (
.O6(p_s0_o15_2),
.O5(),
.I0(a[18]),
.I1(b[0]),
.I2(a[17]),
.I3(b[1]),
.I4(a[16]),
.I5(b[2]));

wire p_s0_o16_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o15_t9_z1_v0 (
.O6(p_s0_o16_0),
.O5(),
.I0(a[18]),
.I1(b[0]),
.I2(a[17]),
.I3(b[1]),
.I4(a[16]),
.I5(b[2]));

wire p_s0_o15_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o15_t9_z0_v1 (
.O6(p_s0_o15_3),
.O5(),
.I0(a[15]),
.I1(b[3]),
.I2(a[14]),
.I3(b[4]),
.I4(a[13]),
.I5(b[5]));

wire p_s0_o16_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o15_t9_z1_v1 (
.O6(p_s0_o16_1),
.O5(),
.I0(a[15]),
.I1(b[3]),
.I2(a[14]),
.I3(b[4]),
.I4(a[13]),
.I5(b[5]));

wire p_s0_o15_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o15_t9_z0_v2 (
.O6(p_s0_o15_4),
.O5(),
.I0(a[12]),
.I1(b[6]),
.I2(a[11]),
.I3(b[7]),
.I4(a[10]),
.I5(b[8]));

wire p_s0_o16_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o15_t9_z1_v2 (
.O6(p_s0_o16_2),
.O5(),
.I0(a[12]),
.I1(b[6]),
.I2(a[11]),
.I3(b[7]),
.I4(a[10]),
.I5(b[8]));

/////////STEP0----ORDER16////////////

wire p_s0_o16_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o16_t10_z0_v0 (
.O6(p_s0_o16_3),
.O5(),
.I0(a[19]),
.I1(b[0]),
.I2(a[18]),
.I3(b[1]),
.I4(a[17]),
.I5(b[2]));

wire p_s0_o17_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o16_t10_z1_v0 (
.O6(p_s0_o17_0),
.O5(),
.I0(a[19]),
.I1(b[0]),
.I2(a[18]),
.I3(b[1]),
.I4(a[17]),
.I5(b[2]));

wire p_s0_o16_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o16_t10_z0_v1 (
.O6(p_s0_o16_4),
.O5(),
.I0(a[16]),
.I1(b[3]),
.I2(a[15]),
.I3(b[4]),
.I4(a[14]),
.I5(b[5]));

wire p_s0_o17_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o16_t10_z1_v1 (
.O6(p_s0_o17_1),
.O5(),
.I0(a[16]),
.I1(b[3]),
.I2(a[15]),
.I3(b[4]),
.I4(a[14]),
.I5(b[5]));

wire p_s0_o16_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o16_t10_z0_v2 (
.O6(p_s0_o16_5),
.O5(),
.I0(a[13]),
.I1(b[6]),
.I2(a[12]),
.I3(b[7]),
.I4(a[11]),
.I5(b[8]));

wire p_s0_o17_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o16_t10_z1_v2 (
.O6(p_s0_o17_2),
.O5(),
.I0(a[13]),
.I1(b[6]),
.I2(a[12]),
.I3(b[7]),
.I4(a[11]),
.I5(b[8]));

/////////STEP0----ORDER17////////////

wire p_s0_o17_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o17_t11_z0_v0 (
.O6(p_s0_o17_3),
.O5(),
.I0(a[20]),
.I1(b[0]),
.I2(a[19]),
.I3(b[1]),
.I4(a[18]),
.I5(b[2]));

wire p_s0_o18_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o17_t11_z1_v0 (
.O6(p_s0_o18_0),
.O5(),
.I0(a[20]),
.I1(b[0]),
.I2(a[19]),
.I3(b[1]),
.I4(a[18]),
.I5(b[2]));

wire p_s0_o17_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o17_t11_z0_v1 (
.O6(p_s0_o17_4),
.O5(),
.I0(a[17]),
.I1(b[3]),
.I2(a[16]),
.I3(b[4]),
.I4(a[15]),
.I5(b[5]));

wire p_s0_o18_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o17_t11_z1_v1 (
.O6(p_s0_o18_1),
.O5(),
.I0(a[17]),
.I1(b[3]),
.I2(a[16]),
.I3(b[4]),
.I4(a[15]),
.I5(b[5]));

wire p_s0_o17_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o17_t11_z0_v2 (
.O6(p_s0_o17_5),
.O5(),
.I0(a[14]),
.I1(b[6]),
.I2(a[13]),
.I3(b[7]),
.I4(a[12]),
.I5(b[8]));

wire p_s0_o18_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o17_t11_z1_v2 (
.O6(p_s0_o18_2),
.O5(),
.I0(a[14]),
.I1(b[6]),
.I2(a[13]),
.I3(b[7]),
.I4(a[12]),
.I5(b[8]));

/////////STEP0----ORDER18////////////

wire p_s0_o18_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o18_t12_z0_v0 (
.O6(p_s0_o18_3),
.O5(),
.I0(a[21]),
.I1(b[0]),
.I2(a[20]),
.I3(b[1]),
.I4(a[19]),
.I5(b[2]));

wire p_s0_o19_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o18_t12_z1_v0 (
.O6(p_s0_o19_0),
.O5(),
.I0(a[21]),
.I1(b[0]),
.I2(a[20]),
.I3(b[1]),
.I4(a[19]),
.I5(b[2]));

wire p_s0_o18_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o18_t12_z0_v1 (
.O6(p_s0_o18_4),
.O5(),
.I0(a[18]),
.I1(b[3]),
.I2(a[17]),
.I3(b[4]),
.I4(a[16]),
.I5(b[5]));

wire p_s0_o19_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o18_t12_z1_v1 (
.O6(p_s0_o19_1),
.O5(),
.I0(a[18]),
.I1(b[3]),
.I2(a[17]),
.I3(b[4]),
.I4(a[16]),
.I5(b[5]));

wire p_s0_o18_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o18_t12_z0_v2 (
.O6(p_s0_o18_5),
.O5(),
.I0(a[15]),
.I1(b[6]),
.I2(a[14]),
.I3(b[7]),
.I4(a[13]),
.I5(b[8]));

wire p_s0_o19_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o18_t12_z1_v2 (
.O6(p_s0_o19_2),
.O5(),
.I0(a[15]),
.I1(b[6]),
.I2(a[14]),
.I3(b[7]),
.I4(a[13]),
.I5(b[8]));

wire p_s0_o18_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o18_t12_z0_v3 (
.O6(p_s0_o18_6),
.O5(),
.I0(a[12]),
.I1(b[9]),
.I2(a[11]),
.I3(b[10]),
.I4(a[10]),
.I5(b[11]));

wire p_s0_o19_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o18_t12_z1_v3 (
.O6(p_s0_o19_3),
.O5(),
.I0(a[12]),
.I1(b[9]),
.I2(a[11]),
.I3(b[10]),
.I4(a[10]),
.I5(b[11]));

/////////STEP0----ORDER19////////////

wire p_s0_o19_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o19_t13_z0_v0 (
.O6(p_s0_o19_4),
.O5(),
.I0(a[22]),
.I1(b[0]),
.I2(a[21]),
.I3(b[1]),
.I4(a[20]),
.I5(b[2]));

wire p_s0_o20_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o19_t13_z1_v0 (
.O6(p_s0_o20_0),
.O5(),
.I0(a[22]),
.I1(b[0]),
.I2(a[21]),
.I3(b[1]),
.I4(a[20]),
.I5(b[2]));

wire p_s0_o19_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o19_t13_z0_v1 (
.O6(p_s0_o19_5),
.O5(),
.I0(a[19]),
.I1(b[3]),
.I2(a[18]),
.I3(b[4]),
.I4(a[17]),
.I5(b[5]));

wire p_s0_o20_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o19_t13_z1_v1 (
.O6(p_s0_o20_1),
.O5(),
.I0(a[19]),
.I1(b[3]),
.I2(a[18]),
.I3(b[4]),
.I4(a[17]),
.I5(b[5]));

wire p_s0_o19_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o19_t13_z0_v2 (
.O6(p_s0_o19_6),
.O5(),
.I0(a[16]),
.I1(b[6]),
.I2(a[15]),
.I3(b[7]),
.I4(a[14]),
.I5(b[8]));

wire p_s0_o20_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o19_t13_z1_v2 (
.O6(p_s0_o20_2),
.O5(),
.I0(a[16]),
.I1(b[6]),
.I2(a[15]),
.I3(b[7]),
.I4(a[14]),
.I5(b[8]));

/////////STEP0----ORDER20////////////

wire p_s0_o20_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o20_t14_z0_v0 (
.O6(p_s0_o20_3),
.O5(),
.I0(a[23]),
.I1(b[0]),
.I2(a[22]),
.I3(b[1]),
.I4(a[21]),
.I5(b[2]));

wire p_s0_o21_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o20_t14_z1_v0 (
.O6(p_s0_o21_0),
.O5(),
.I0(a[23]),
.I1(b[0]),
.I2(a[22]),
.I3(b[1]),
.I4(a[21]),
.I5(b[2]));

wire p_s0_o20_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o20_t14_z0_v1 (
.O6(p_s0_o20_4),
.O5(),
.I0(a[20]),
.I1(b[3]),
.I2(a[19]),
.I3(b[4]),
.I4(a[18]),
.I5(b[5]));

wire p_s0_o21_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o20_t14_z1_v1 (
.O6(p_s0_o21_1),
.O5(),
.I0(a[20]),
.I1(b[3]),
.I2(a[19]),
.I3(b[4]),
.I4(a[18]),
.I5(b[5]));

wire p_s0_o20_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o20_t14_z0_v2 (
.O6(p_s0_o20_5),
.O5(),
.I0(a[17]),
.I1(b[6]),
.I2(a[16]),
.I3(b[7]),
.I4(a[15]),
.I5(b[8]));

wire p_s0_o21_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o20_t14_z1_v2 (
.O6(p_s0_o21_2),
.O5(),
.I0(a[17]),
.I1(b[6]),
.I2(a[16]),
.I3(b[7]),
.I4(a[15]),
.I5(b[8]));

wire p_s0_o20_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o20_t14_z0_v3 (
.O6(p_s0_o20_6),
.O5(),
.I0(a[14]),
.I1(b[9]),
.I2(a[13]),
.I3(b[10]),
.I4(a[12]),
.I5(b[11]));

wire p_s0_o21_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o20_t14_z1_v3 (
.O6(p_s0_o21_3),
.O5(),
.I0(a[14]),
.I1(b[9]),
.I2(a[13]),
.I3(b[10]),
.I4(a[12]),
.I5(b[11]));

wire p_s0_o20_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o20_t14_z0_v4 (
.O6(p_s0_o20_7),
.O5(),
.I0(a[11]),
.I1(b[12]),
.I2(a[10]),
.I3(b[13]),
.I4(a[9]),
.I5(b[14]));

wire p_s0_o21_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o20_t14_z1_v4 (
.O6(p_s0_o21_4),
.O5(),
.I0(a[11]),
.I1(b[12]),
.I2(a[10]),
.I3(b[13]),
.I4(a[9]),
.I5(b[14]));

wire p_s0_o20_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o20_t14_z0_v5 (
.O6(p_s0_o20_8),
.O5(),
.I0(a[8]),
.I1(b[15]),
.I2(a[7]),
.I3(b[16]),
.I4(a[6]),
.I5(b[17]));

wire p_s0_o21_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o20_t14_z1_v5 (
.O6(p_s0_o21_5),
.O5(),
.I0(a[8]),
.I1(b[15]),
.I2(a[7]),
.I3(b[16]),
.I4(a[6]),
.I5(b[17]));

/////////STEP0----ORDER21////////////

wire p_s0_o21_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o21_t15_z0_v0 (
.O6(p_s0_o21_6),
.O5(),
.I0(a[24]),
.I1(b[0]),
.I2(a[23]),
.I3(b[1]),
.I4(a[22]),
.I5(b[2]));

wire p_s0_o22_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o21_t15_z1_v0 (
.O6(p_s0_o22_0),
.O5(),
.I0(a[24]),
.I1(b[0]),
.I2(a[23]),
.I3(b[1]),
.I4(a[22]),
.I5(b[2]));

wire p_s0_o21_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o21_t15_z0_v1 (
.O6(p_s0_o21_7),
.O5(),
.I0(a[21]),
.I1(b[3]),
.I2(a[20]),
.I3(b[4]),
.I4(a[19]),
.I5(b[5]));

wire p_s0_o22_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o21_t15_z1_v1 (
.O6(p_s0_o22_1),
.O5(),
.I0(a[21]),
.I1(b[3]),
.I2(a[20]),
.I3(b[4]),
.I4(a[19]),
.I5(b[5]));

wire p_s0_o21_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o21_t15_z0_v2 (
.O6(p_s0_o21_8),
.O5(),
.I0(a[18]),
.I1(b[6]),
.I2(a[17]),
.I3(b[7]),
.I4(a[16]),
.I5(b[8]));

wire p_s0_o22_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o21_t15_z1_v2 (
.O6(p_s0_o22_2),
.O5(),
.I0(a[18]),
.I1(b[6]),
.I2(a[17]),
.I3(b[7]),
.I4(a[16]),
.I5(b[8]));

/////////STEP0----ORDER22////////////

wire p_s0_o22_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t16_z0_v0 (
.O6(p_s0_o22_3),
.O5(),
.I0(a[25]),
.I1(b[0]),
.I2(a[24]),
.I3(b[1]),
.I4(a[23]),
.I5(b[2]));

wire p_s0_o23_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t16_z1_v0 (
.O6(p_s0_o23_0),
.O5(),
.I0(a[25]),
.I1(b[0]),
.I2(a[24]),
.I3(b[1]),
.I4(a[23]),
.I5(b[2]));

wire p_s0_o22_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t16_z0_v1 (
.O6(p_s0_o22_4),
.O5(),
.I0(a[22]),
.I1(b[3]),
.I2(a[21]),
.I3(b[4]),
.I4(a[20]),
.I5(b[5]));

wire p_s0_o23_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t16_z1_v1 (
.O6(p_s0_o23_1),
.O5(),
.I0(a[22]),
.I1(b[3]),
.I2(a[21]),
.I3(b[4]),
.I4(a[20]),
.I5(b[5]));

wire p_s0_o22_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t16_z0_v2 (
.O6(p_s0_o22_5),
.O5(),
.I0(a[19]),
.I1(b[6]),
.I2(a[18]),
.I3(b[7]),
.I4(a[17]),
.I5(b[8]));

wire p_s0_o23_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t16_z1_v2 (
.O6(p_s0_o23_2),
.O5(),
.I0(a[19]),
.I1(b[6]),
.I2(a[18]),
.I3(b[7]),
.I4(a[17]),
.I5(b[8]));

wire p_s0_o22_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t16_z0_v3 (
.O6(p_s0_o22_6),
.O5(),
.I0(a[16]),
.I1(b[9]),
.I2(a[15]),
.I3(b[10]),
.I4(a[14]),
.I5(b[11]));

wire p_s0_o23_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t16_z1_v3 (
.O6(p_s0_o23_3),
.O5(),
.I0(a[16]),
.I1(b[9]),
.I2(a[15]),
.I3(b[10]),
.I4(a[14]),
.I5(b[11]));

wire p_s0_o22_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t16_z0_v4 (
.O6(p_s0_o22_7),
.O5(),
.I0(a[13]),
.I1(b[12]),
.I2(a[12]),
.I3(b[13]),
.I4(a[11]),
.I5(b[14]));

wire p_s0_o23_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t16_z1_v4 (
.O6(p_s0_o23_4),
.O5(),
.I0(a[13]),
.I1(b[12]),
.I2(a[12]),
.I3(b[13]),
.I4(a[11]),
.I5(b[14]));

wire p_s0_o22_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t16_z0_v5 (
.O6(p_s0_o22_8),
.O5(),
.I0(a[10]),
.I1(b[15]),
.I2(a[9]),
.I3(b[16]),
.I4(a[8]),
.I5(b[17]));

wire p_s0_o23_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t16_z1_v5 (
.O6(p_s0_o23_5),
.O5(),
.I0(a[10]),
.I1(b[15]),
.I2(a[9]),
.I3(b[16]),
.I4(a[8]),
.I5(b[17]));

wire p_s0_o22_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t16_z0_v6 (
.O6(p_s0_o22_9),
.O5(),
.I0(a[7]),
.I1(b[18]),
.I2(a[6]),
.I3(b[19]),
.I4(a[5]),
.I5(b[20]));

wire p_s0_o23_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t16_z1_v6 (
.O6(p_s0_o23_6),
.O5(),
.I0(a[7]),
.I1(b[18]),
.I2(a[6]),
.I3(b[19]),
.I4(a[5]),
.I5(b[20]));

wire p_s0_o22_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t16_z0_v7 (
.O6(p_s0_o22_10),
.O5(),
.I0(a[4]),
.I1(b[21]),
.I2(a[3]),
.I3(b[22]),
.I4(a[2]),
.I5(b[23]));

wire p_s0_o23_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t16_z1_v7 (
.O6(p_s0_o23_7),
.O5(),
.I0(a[4]),
.I1(b[21]),
.I2(a[3]),
.I3(b[22]),
.I4(a[2]),
.I5(b[23]));

/////////STEP0----ORDER23////////////

wire p_s0_o23_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o23_t17_z0_v0 (
.O6(p_s0_o23_8),
.O5(),
.I0(a[26]),
.I1(b[0]),
.I2(a[25]),
.I3(b[1]),
.I4(a[24]),
.I5(b[2]));

wire p_s0_o24_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o23_t17_z1_v0 (
.O6(p_s0_o24_0),
.O5(),
.I0(a[26]),
.I1(b[0]),
.I2(a[25]),
.I3(b[1]),
.I4(a[24]),
.I5(b[2]));

wire p_s0_o23_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o23_t17_z0_v1 (
.O6(p_s0_o23_9),
.O5(),
.I0(a[23]),
.I1(b[3]),
.I2(a[22]),
.I3(b[4]),
.I4(a[21]),
.I5(b[5]));

wire p_s0_o24_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o23_t17_z1_v1 (
.O6(p_s0_o24_1),
.O5(),
.I0(a[23]),
.I1(b[3]),
.I2(a[22]),
.I3(b[4]),
.I4(a[21]),
.I5(b[5]));

wire p_s0_o23_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o23_t17_z0_v2 (
.O6(p_s0_o23_10),
.O5(),
.I0(a[20]),
.I1(b[6]),
.I2(a[19]),
.I3(b[7]),
.I4(a[18]),
.I5(b[8]));

wire p_s0_o24_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o23_t17_z1_v2 (
.O6(p_s0_o24_2),
.O5(),
.I0(a[20]),
.I1(b[6]),
.I2(a[19]),
.I3(b[7]),
.I4(a[18]),
.I5(b[8]));

wire p_s0_o23_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o23_t17_z0_v3 (
.O6(p_s0_o23_11),
.O5(),
.I0(a[17]),
.I1(b[9]),
.I2(a[16]),
.I3(b[10]),
.I4(a[15]),
.I5(b[11]));

wire p_s0_o24_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o23_t17_z1_v3 (
.O6(p_s0_o24_3),
.O5(),
.I0(a[17]),
.I1(b[9]),
.I2(a[16]),
.I3(b[10]),
.I4(a[15]),
.I5(b[11]));

wire p_s0_o23_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o23_t17_z0_v4 (
.O6(p_s0_o23_12),
.O5(),
.I0(a[14]),
.I1(b[12]),
.I2(a[13]),
.I3(b[13]),
.I4(a[12]),
.I5(b[14]));

wire p_s0_o24_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o23_t17_z1_v4 (
.O6(p_s0_o24_4),
.O5(),
.I0(a[14]),
.I1(b[12]),
.I2(a[13]),
.I3(b[13]),
.I4(a[12]),
.I5(b[14]));

/////////STEP0----ORDER24////////////

wire p_s0_o24_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v0 (
.O6(p_s0_o24_5),
.O5(),
.I0(a[27]),
.I1(b[0]),
.I2(a[26]),
.I3(b[1]),
.I4(a[25]),
.I5(b[2]));

wire p_s0_o25_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v0 (
.O6(p_s0_o25_0),
.O5(),
.I0(a[27]),
.I1(b[0]),
.I2(a[26]),
.I3(b[1]),
.I4(a[25]),
.I5(b[2]));

wire p_s0_o24_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v1 (
.O6(p_s0_o24_6),
.O5(),
.I0(a[24]),
.I1(b[3]),
.I2(a[23]),
.I3(b[4]),
.I4(a[22]),
.I5(b[5]));

wire p_s0_o25_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v1 (
.O6(p_s0_o25_1),
.O5(),
.I0(a[24]),
.I1(b[3]),
.I2(a[23]),
.I3(b[4]),
.I4(a[22]),
.I5(b[5]));

wire p_s0_o24_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v2 (
.O6(p_s0_o24_7),
.O5(),
.I0(a[21]),
.I1(b[6]),
.I2(a[20]),
.I3(b[7]),
.I4(a[19]),
.I5(b[8]));

wire p_s0_o25_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v2 (
.O6(p_s0_o25_2),
.O5(),
.I0(a[21]),
.I1(b[6]),
.I2(a[20]),
.I3(b[7]),
.I4(a[19]),
.I5(b[8]));

wire p_s0_o24_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v3 (
.O6(p_s0_o24_8),
.O5(),
.I0(a[18]),
.I1(b[9]),
.I2(a[17]),
.I3(b[10]),
.I4(a[16]),
.I5(b[11]));

wire p_s0_o25_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v3 (
.O6(p_s0_o25_3),
.O5(),
.I0(a[18]),
.I1(b[9]),
.I2(a[17]),
.I3(b[10]),
.I4(a[16]),
.I5(b[11]));

wire p_s0_o24_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v4 (
.O6(p_s0_o24_9),
.O5(),
.I0(a[15]),
.I1(b[12]),
.I2(a[14]),
.I3(b[13]),
.I4(a[13]),
.I5(b[14]));

wire p_s0_o25_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v4 (
.O6(p_s0_o25_4),
.O5(),
.I0(a[15]),
.I1(b[12]),
.I2(a[14]),
.I3(b[13]),
.I4(a[13]),
.I5(b[14]));

wire p_s0_o24_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v5 (
.O6(p_s0_o24_10),
.O5(),
.I0(a[12]),
.I1(b[15]),
.I2(a[11]),
.I3(b[16]),
.I4(a[10]),
.I5(b[17]));

wire p_s0_o25_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v5 (
.O6(p_s0_o25_5),
.O5(),
.I0(a[12]),
.I1(b[15]),
.I2(a[11]),
.I3(b[16]),
.I4(a[10]),
.I5(b[17]));

wire p_s0_o24_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v6 (
.O6(p_s0_o24_11),
.O5(),
.I0(a[9]),
.I1(b[18]),
.I2(a[8]),
.I3(b[19]),
.I4(a[7]),
.I5(b[20]));

wire p_s0_o25_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v6 (
.O6(p_s0_o25_6),
.O5(),
.I0(a[9]),
.I1(b[18]),
.I2(a[8]),
.I3(b[19]),
.I4(a[7]),
.I5(b[20]));

wire p_s0_o24_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v7 (
.O6(p_s0_o24_12),
.O5(),
.I0(a[6]),
.I1(b[21]),
.I2(a[5]),
.I3(b[22]),
.I4(a[4]),
.I5(b[23]));

wire p_s0_o25_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v7 (
.O6(p_s0_o25_7),
.O5(),
.I0(a[6]),
.I1(b[21]),
.I2(a[5]),
.I3(b[22]),
.I4(a[4]),
.I5(b[23]));

wire p_s0_o24_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o24_t18_z0_v8 (
.O6(p_s0_o24_13),
.O5(),
.I0(a[3]),
.I1(b[24]),
.I2(a[2]),
.I3(b[25]),
.I4(a[1]),
.I5(b[26]));

wire p_s0_o25_8;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o24_t18_z1_v8 (
.O6(p_s0_o25_8),
.O5(),
.I0(a[3]),
.I1(b[24]),
.I2(a[2]),
.I3(b[25]),
.I4(a[1]),
.I5(b[26]));

/////////STEP0----ORDER25////////////

wire p_s0_o25_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o25_t19_z0_v0 (
.O6(p_s0_o25_9),
.O5(),
.I0(a[28]),
.I1(b[0]),
.I2(a[27]),
.I3(b[1]),
.I4(a[26]),
.I5(b[2]));

wire p_s0_o26_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o25_t19_z1_v0 (
.O6(p_s0_o26_0),
.O5(),
.I0(a[28]),
.I1(b[0]),
.I2(a[27]),
.I3(b[1]),
.I4(a[26]),
.I5(b[2]));

wire p_s0_o25_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o25_t19_z0_v1 (
.O6(p_s0_o25_10),
.O5(),
.I0(a[25]),
.I1(b[3]),
.I2(a[24]),
.I3(b[4]),
.I4(a[23]),
.I5(b[5]));

wire p_s0_o26_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o25_t19_z1_v1 (
.O6(p_s0_o26_1),
.O5(),
.I0(a[25]),
.I1(b[3]),
.I2(a[24]),
.I3(b[4]),
.I4(a[23]),
.I5(b[5]));

wire p_s0_o25_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o25_t19_z0_v2 (
.O6(p_s0_o25_11),
.O5(),
.I0(a[22]),
.I1(b[6]),
.I2(a[21]),
.I3(b[7]),
.I4(a[20]),
.I5(b[8]));

wire p_s0_o26_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o25_t19_z1_v2 (
.O6(p_s0_o26_2),
.O5(),
.I0(a[22]),
.I1(b[6]),
.I2(a[21]),
.I3(b[7]),
.I4(a[20]),
.I5(b[8]));

/////////STEP0----ORDER26////////////

wire p_s0_o26_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v0 (
.O6(p_s0_o26_3),
.O5(),
.I0(a[29]),
.I1(b[0]),
.I2(a[28]),
.I3(b[1]),
.I4(a[27]),
.I5(b[2]));

wire p_s0_o27_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v0 (
.O6(p_s0_o27_0),
.O5(),
.I0(a[29]),
.I1(b[0]),
.I2(a[28]),
.I3(b[1]),
.I4(a[27]),
.I5(b[2]));

wire p_s0_o26_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v1 (
.O6(p_s0_o26_4),
.O5(),
.I0(a[26]),
.I1(b[3]),
.I2(a[25]),
.I3(b[4]),
.I4(a[24]),
.I5(b[5]));

wire p_s0_o27_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v1 (
.O6(p_s0_o27_1),
.O5(),
.I0(a[26]),
.I1(b[3]),
.I2(a[25]),
.I3(b[4]),
.I4(a[24]),
.I5(b[5]));

wire p_s0_o26_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v2 (
.O6(p_s0_o26_5),
.O5(),
.I0(a[23]),
.I1(b[6]),
.I2(a[22]),
.I3(b[7]),
.I4(a[21]),
.I5(b[8]));

wire p_s0_o27_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v2 (
.O6(p_s0_o27_2),
.O5(),
.I0(a[23]),
.I1(b[6]),
.I2(a[22]),
.I3(b[7]),
.I4(a[21]),
.I5(b[8]));

wire p_s0_o26_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v3 (
.O6(p_s0_o26_6),
.O5(),
.I0(a[20]),
.I1(b[9]),
.I2(a[19]),
.I3(b[10]),
.I4(a[18]),
.I5(b[11]));

wire p_s0_o27_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v3 (
.O6(p_s0_o27_3),
.O5(),
.I0(a[20]),
.I1(b[9]),
.I2(a[19]),
.I3(b[10]),
.I4(a[18]),
.I5(b[11]));

wire p_s0_o26_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v4 (
.O6(p_s0_o26_7),
.O5(),
.I0(a[17]),
.I1(b[12]),
.I2(a[16]),
.I3(b[13]),
.I4(a[15]),
.I5(b[14]));

wire p_s0_o27_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v4 (
.O6(p_s0_o27_4),
.O5(),
.I0(a[17]),
.I1(b[12]),
.I2(a[16]),
.I3(b[13]),
.I4(a[15]),
.I5(b[14]));

wire p_s0_o26_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v5 (
.O6(p_s0_o26_8),
.O5(),
.I0(a[14]),
.I1(b[15]),
.I2(a[13]),
.I3(b[16]),
.I4(a[12]),
.I5(b[17]));

wire p_s0_o27_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v5 (
.O6(p_s0_o27_5),
.O5(),
.I0(a[14]),
.I1(b[15]),
.I2(a[13]),
.I3(b[16]),
.I4(a[12]),
.I5(b[17]));

wire p_s0_o26_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v6 (
.O6(p_s0_o26_9),
.O5(),
.I0(a[11]),
.I1(b[18]),
.I2(a[10]),
.I3(b[19]),
.I4(a[9]),
.I5(b[20]));

wire p_s0_o27_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v6 (
.O6(p_s0_o27_6),
.O5(),
.I0(a[11]),
.I1(b[18]),
.I2(a[10]),
.I3(b[19]),
.I4(a[9]),
.I5(b[20]));

wire p_s0_o26_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v7 (
.O6(p_s0_o26_10),
.O5(),
.I0(a[8]),
.I1(b[21]),
.I2(a[7]),
.I3(b[22]),
.I4(a[6]),
.I5(b[23]));

wire p_s0_o27_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v7 (
.O6(p_s0_o27_7),
.O5(),
.I0(a[8]),
.I1(b[21]),
.I2(a[7]),
.I3(b[22]),
.I4(a[6]),
.I5(b[23]));

wire p_s0_o26_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v8 (
.O6(p_s0_o26_11),
.O5(),
.I0(a[5]),
.I1(b[24]),
.I2(a[4]),
.I3(b[25]),
.I4(a[3]),
.I5(b[26]));

wire p_s0_o27_8;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v8 (
.O6(p_s0_o27_8),
.O5(),
.I0(a[5]),
.I1(b[24]),
.I2(a[4]),
.I3(b[25]),
.I4(a[3]),
.I5(b[26]));

wire p_s0_o26_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o26_t20_z0_v9 (
.O6(p_s0_o26_12),
.O5(),
.I0(a[2]),
.I1(b[27]),
.I2(a[1]),
.I3(b[28]),
.I4(a[0]),
.I5(b[29]));

wire p_s0_o27_9;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o26_t20_z1_v9 (
.O6(p_s0_o27_9),
.O5(),
.I0(a[2]),
.I1(b[27]),
.I2(a[1]),
.I3(b[28]),
.I4(a[0]),
.I5(b[29]));

/////////STEP0----ORDER27////////////

wire p_s0_o27_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v0 (
.O6(p_s0_o27_10),
.O5(),
.I0(a[30]),
.I1(b[0]),
.I2(a[29]),
.I3(b[1]),
.I4(a[28]),
.I5(b[2]));

wire p_s0_o28_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v0 (
.O6(p_s0_o28_0),
.O5(),
.I0(a[30]),
.I1(b[0]),
.I2(a[29]),
.I3(b[1]),
.I4(a[28]),
.I5(b[2]));

wire p_s0_o27_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v1 (
.O6(p_s0_o27_11),
.O5(),
.I0(a[27]),
.I1(b[3]),
.I2(a[26]),
.I3(b[4]),
.I4(a[25]),
.I5(b[5]));

wire p_s0_o28_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v1 (
.O6(p_s0_o28_1),
.O5(),
.I0(a[27]),
.I1(b[3]),
.I2(a[26]),
.I3(b[4]),
.I4(a[25]),
.I5(b[5]));

wire p_s0_o27_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v2 (
.O6(p_s0_o27_12),
.O5(),
.I0(a[24]),
.I1(b[6]),
.I2(a[23]),
.I3(b[7]),
.I4(a[22]),
.I5(b[8]));

wire p_s0_o28_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v2 (
.O6(p_s0_o28_2),
.O5(),
.I0(a[24]),
.I1(b[6]),
.I2(a[23]),
.I3(b[7]),
.I4(a[22]),
.I5(b[8]));

wire p_s0_o27_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v3 (
.O6(p_s0_o27_13),
.O5(),
.I0(a[21]),
.I1(b[9]),
.I2(a[20]),
.I3(b[10]),
.I4(a[19]),
.I5(b[11]));

wire p_s0_o28_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v3 (
.O6(p_s0_o28_3),
.O5(),
.I0(a[21]),
.I1(b[9]),
.I2(a[20]),
.I3(b[10]),
.I4(a[19]),
.I5(b[11]));

wire p_s0_o27_14;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v4 (
.O6(p_s0_o27_14),
.O5(),
.I0(a[18]),
.I1(b[12]),
.I2(a[17]),
.I3(b[13]),
.I4(a[16]),
.I5(b[14]));

wire p_s0_o28_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v4 (
.O6(p_s0_o28_4),
.O5(),
.I0(a[18]),
.I1(b[12]),
.I2(a[17]),
.I3(b[13]),
.I4(a[16]),
.I5(b[14]));

wire p_s0_o27_15;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v5 (
.O6(p_s0_o27_15),
.O5(),
.I0(a[15]),
.I1(b[15]),
.I2(a[14]),
.I3(b[16]),
.I4(a[13]),
.I5(b[17]));

wire p_s0_o28_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v5 (
.O6(p_s0_o28_5),
.O5(),
.I0(a[15]),
.I1(b[15]),
.I2(a[14]),
.I3(b[16]),
.I4(a[13]),
.I5(b[17]));

wire p_s0_o27_16;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v6 (
.O6(p_s0_o27_16),
.O5(),
.I0(a[12]),
.I1(b[18]),
.I2(a[11]),
.I3(b[19]),
.I4(a[10]),
.I5(b[20]));

wire p_s0_o28_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v6 (
.O6(p_s0_o28_6),
.O5(),
.I0(a[12]),
.I1(b[18]),
.I2(a[11]),
.I3(b[19]),
.I4(a[10]),
.I5(b[20]));

wire p_s0_o27_17;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v7 (
.O6(p_s0_o27_17),
.O5(),
.I0(a[9]),
.I1(b[21]),
.I2(a[8]),
.I3(b[22]),
.I4(a[7]),
.I5(b[23]));

wire p_s0_o28_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v7 (
.O6(p_s0_o28_7),
.O5(),
.I0(a[9]),
.I1(b[21]),
.I2(a[8]),
.I3(b[22]),
.I4(a[7]),
.I5(b[23]));

wire p_s0_o27_18;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o27_t21_z0_v8 (
.O6(p_s0_o27_18),
.O5(),
.I0(a[6]),
.I1(b[24]),
.I2(a[5]),
.I3(b[25]),
.I4(a[4]),
.I5(b[26]));

wire p_s0_o28_8;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o27_t21_z1_v8 (
.O6(p_s0_o28_8),
.O5(),
.I0(a[6]),
.I1(b[24]),
.I2(a[5]),
.I3(b[25]),
.I4(a[4]),
.I5(b[26]));

/////////STEP0----ORDER28////////////

wire p_s0_o28_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v0 (
.O6(p_s0_o28_9),
.O5(),
.I0(a[31]),
.I1(b[0]),
.I2(a[30]),
.I3(b[1]),
.I4(a[29]),
.I5(b[2]));

wire p_s0_o29_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v0 (
.O6(p_s0_o29_0),
.O5(),
.I0(a[31]),
.I1(b[0]),
.I2(a[30]),
.I3(b[1]),
.I4(a[29]),
.I5(b[2]));

wire p_s0_o28_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v1 (
.O6(p_s0_o28_10),
.O5(),
.I0(a[28]),
.I1(b[3]),
.I2(a[27]),
.I3(b[4]),
.I4(a[26]),
.I5(b[5]));

wire p_s0_o29_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v1 (
.O6(p_s0_o29_1),
.O5(),
.I0(a[28]),
.I1(b[3]),
.I2(a[27]),
.I3(b[4]),
.I4(a[26]),
.I5(b[5]));

wire p_s0_o28_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v2 (
.O6(p_s0_o28_11),
.O5(),
.I0(a[25]),
.I1(b[6]),
.I2(a[24]),
.I3(b[7]),
.I4(a[23]),
.I5(b[8]));

wire p_s0_o29_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v2 (
.O6(p_s0_o29_2),
.O5(),
.I0(a[25]),
.I1(b[6]),
.I2(a[24]),
.I3(b[7]),
.I4(a[23]),
.I5(b[8]));

wire p_s0_o28_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v3 (
.O6(p_s0_o28_12),
.O5(),
.I0(a[22]),
.I1(b[9]),
.I2(a[21]),
.I3(b[10]),
.I4(a[20]),
.I5(b[11]));

wire p_s0_o29_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v3 (
.O6(p_s0_o29_3),
.O5(),
.I0(a[22]),
.I1(b[9]),
.I2(a[21]),
.I3(b[10]),
.I4(a[20]),
.I5(b[11]));

wire p_s0_o28_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v4 (
.O6(p_s0_o28_13),
.O5(),
.I0(a[19]),
.I1(b[12]),
.I2(a[18]),
.I3(b[13]),
.I4(a[17]),
.I5(b[14]));

wire p_s0_o29_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v4 (
.O6(p_s0_o29_4),
.O5(),
.I0(a[19]),
.I1(b[12]),
.I2(a[18]),
.I3(b[13]),
.I4(a[17]),
.I5(b[14]));

wire p_s0_o28_14;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v5 (
.O6(p_s0_o28_14),
.O5(),
.I0(a[16]),
.I1(b[15]),
.I2(a[15]),
.I3(b[16]),
.I4(a[14]),
.I5(b[17]));

wire p_s0_o29_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v5 (
.O6(p_s0_o29_5),
.O5(),
.I0(a[16]),
.I1(b[15]),
.I2(a[15]),
.I3(b[16]),
.I4(a[14]),
.I5(b[17]));

wire p_s0_o28_15;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v6 (
.O6(p_s0_o28_15),
.O5(),
.I0(a[13]),
.I1(b[18]),
.I2(a[12]),
.I3(b[19]),
.I4(a[11]),
.I5(b[20]));

wire p_s0_o29_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v6 (
.O6(p_s0_o29_6),
.O5(),
.I0(a[13]),
.I1(b[18]),
.I2(a[12]),
.I3(b[19]),
.I4(a[11]),
.I5(b[20]));

wire p_s0_o28_16;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v7 (
.O6(p_s0_o28_16),
.O5(),
.I0(a[10]),
.I1(b[21]),
.I2(a[9]),
.I3(b[22]),
.I4(a[8]),
.I5(b[23]));

wire p_s0_o29_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v7 (
.O6(p_s0_o29_7),
.O5(),
.I0(a[10]),
.I1(b[21]),
.I2(a[9]),
.I3(b[22]),
.I4(a[8]),
.I5(b[23]));

wire p_s0_o28_17;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v8 (
.O6(p_s0_o28_17),
.O5(),
.I0(a[7]),
.I1(b[24]),
.I2(a[6]),
.I3(b[25]),
.I4(a[5]),
.I5(b[26]));

wire p_s0_o29_8;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v8 (
.O6(p_s0_o29_8),
.O5(),
.I0(a[7]),
.I1(b[24]),
.I2(a[6]),
.I3(b[25]),
.I4(a[5]),
.I5(b[26]));

wire p_s0_o28_18;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o28_t22_z0_v9 (
.O6(p_s0_o28_18),
.O5(),
.I0(a[4]),
.I1(b[27]),
.I2(a[3]),
.I3(b[28]),
.I4(a[2]),
.I5(b[29]));

wire p_s0_o29_9;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o28_t22_z1_v9 (
.O6(p_s0_o29_9),
.O5(),
.I0(a[4]),
.I1(b[27]),
.I2(a[3]),
.I3(b[28]),
.I4(a[2]),
.I5(b[29]));

/////////STEP0----ORDER29////////////

wire p_s0_o29_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v0 (
.O6(p_s0_o29_10),
.O5(),
.I0(a[31]),
.I1(b[1]),
.I2(a[30]),
.I3(b[2]),
.I4(a[29]),
.I5(b[3]));

wire p_s0_o30_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v0 (
.O6(p_s0_o30_0),
.O5(),
.I0(a[31]),
.I1(b[1]),
.I2(a[30]),
.I3(b[2]),
.I4(a[29]),
.I5(b[3]));

wire p_s0_o29_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v1 (
.O6(p_s0_o29_11),
.O5(),
.I0(a[28]),
.I1(b[4]),
.I2(a[27]),
.I3(b[5]),
.I4(a[26]),
.I5(b[6]));

wire p_s0_o30_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v1 (
.O6(p_s0_o30_1),
.O5(),
.I0(a[28]),
.I1(b[4]),
.I2(a[27]),
.I3(b[5]),
.I4(a[26]),
.I5(b[6]));

wire p_s0_o29_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v2 (
.O6(p_s0_o29_12),
.O5(),
.I0(a[25]),
.I1(b[7]),
.I2(a[24]),
.I3(b[8]),
.I4(a[23]),
.I5(b[9]));

wire p_s0_o30_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v2 (
.O6(p_s0_o30_2),
.O5(),
.I0(a[25]),
.I1(b[7]),
.I2(a[24]),
.I3(b[8]),
.I4(a[23]),
.I5(b[9]));

wire p_s0_o29_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v3 (
.O6(p_s0_o29_13),
.O5(),
.I0(a[22]),
.I1(b[10]),
.I2(a[21]),
.I3(b[11]),
.I4(a[20]),
.I5(b[12]));

wire p_s0_o30_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v3 (
.O6(p_s0_o30_3),
.O5(),
.I0(a[22]),
.I1(b[10]),
.I2(a[21]),
.I3(b[11]),
.I4(a[20]),
.I5(b[12]));

wire p_s0_o29_14;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v4 (
.O6(p_s0_o29_14),
.O5(),
.I0(a[19]),
.I1(b[13]),
.I2(a[18]),
.I3(b[14]),
.I4(a[17]),
.I5(b[15]));

wire p_s0_o30_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v4 (
.O6(p_s0_o30_4),
.O5(),
.I0(a[19]),
.I1(b[13]),
.I2(a[18]),
.I3(b[14]),
.I4(a[17]),
.I5(b[15]));

wire p_s0_o29_15;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v5 (
.O6(p_s0_o29_15),
.O5(),
.I0(a[16]),
.I1(b[16]),
.I2(a[15]),
.I3(b[17]),
.I4(a[14]),
.I5(b[18]));

wire p_s0_o30_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v5 (
.O6(p_s0_o30_5),
.O5(),
.I0(a[16]),
.I1(b[16]),
.I2(a[15]),
.I3(b[17]),
.I4(a[14]),
.I5(b[18]));

wire p_s0_o29_16;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v6 (
.O6(p_s0_o29_16),
.O5(),
.I0(a[13]),
.I1(b[19]),
.I2(a[12]),
.I3(b[20]),
.I4(a[11]),
.I5(b[21]));

wire p_s0_o30_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v6 (
.O6(p_s0_o30_6),
.O5(),
.I0(a[13]),
.I1(b[19]),
.I2(a[12]),
.I3(b[20]),
.I4(a[11]),
.I5(b[21]));

wire p_s0_o29_17;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v7 (
.O6(p_s0_o29_17),
.O5(),
.I0(a[10]),
.I1(b[22]),
.I2(a[9]),
.I3(b[23]),
.I4(a[8]),
.I5(b[24]));

wire p_s0_o30_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v7 (
.O6(p_s0_o30_7),
.O5(),
.I0(a[10]),
.I1(b[22]),
.I2(a[9]),
.I3(b[23]),
.I4(a[8]),
.I5(b[24]));

wire p_s0_o29_18;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v8 (
.O6(p_s0_o29_18),
.O5(),
.I0(a[7]),
.I1(b[25]),
.I2(a[6]),
.I3(b[26]),
.I4(a[5]),
.I5(b[27]));

wire p_s0_o30_8;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v8 (
.O6(p_s0_o30_8),
.O5(),
.I0(a[7]),
.I1(b[25]),
.I2(a[6]),
.I3(b[26]),
.I4(a[5]),
.I5(b[27]));

wire p_s0_o29_19;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o29_t23_z0_v9 (
.O6(p_s0_o29_19),
.O5(),
.I0(a[4]),
.I1(b[28]),
.I2(a[3]),
.I3(b[29]),
.I4(a[2]),
.I5(b[30]));

wire p_s0_o30_9;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o29_t23_z1_v9 (
.O6(p_s0_o30_9),
.O5(),
.I0(a[4]),
.I1(b[28]),
.I2(a[3]),
.I3(b[29]),
.I4(a[2]),
.I5(b[30]));

/////////STEP0----ORDER30////////////

wire p_s0_o30_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v0 (
.O6(p_s0_o30_10),
.O5(),
.I0(a[31]),
.I1(b[2]),
.I2(a[30]),
.I3(b[3]),
.I4(a[29]),
.I5(b[4]));

wire p_s0_o31_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v0 (
.O6(p_s0_o31_0),
.O5(),
.I0(a[31]),
.I1(b[2]),
.I2(a[30]),
.I3(b[3]),
.I4(a[29]),
.I5(b[4]));

wire p_s0_o30_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v1 (
.O6(p_s0_o30_11),
.O5(),
.I0(a[28]),
.I1(b[5]),
.I2(a[27]),
.I3(b[6]),
.I4(a[26]),
.I5(b[7]));

wire p_s0_o31_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v1 (
.O6(p_s0_o31_1),
.O5(),
.I0(a[28]),
.I1(b[5]),
.I2(a[27]),
.I3(b[6]),
.I4(a[26]),
.I5(b[7]));

wire p_s0_o30_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v2 (
.O6(p_s0_o30_12),
.O5(),
.I0(a[25]),
.I1(b[8]),
.I2(a[24]),
.I3(b[9]),
.I4(a[23]),
.I5(b[10]));

wire p_s0_o31_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v2 (
.O6(p_s0_o31_2),
.O5(),
.I0(a[25]),
.I1(b[8]),
.I2(a[24]),
.I3(b[9]),
.I4(a[23]),
.I5(b[10]));

wire p_s0_o30_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v3 (
.O6(p_s0_o30_13),
.O5(),
.I0(a[22]),
.I1(b[11]),
.I2(a[21]),
.I3(b[12]),
.I4(a[20]),
.I5(b[13]));

wire p_s0_o31_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v3 (
.O6(p_s0_o31_3),
.O5(),
.I0(a[22]),
.I1(b[11]),
.I2(a[21]),
.I3(b[12]),
.I4(a[20]),
.I5(b[13]));

wire p_s0_o30_14;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v4 (
.O6(p_s0_o30_14),
.O5(),
.I0(a[19]),
.I1(b[14]),
.I2(a[18]),
.I3(b[15]),
.I4(a[17]),
.I5(b[16]));

wire p_s0_o31_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v4 (
.O6(p_s0_o31_4),
.O5(),
.I0(a[19]),
.I1(b[14]),
.I2(a[18]),
.I3(b[15]),
.I4(a[17]),
.I5(b[16]));

wire p_s0_o30_15;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v5 (
.O6(p_s0_o30_15),
.O5(),
.I0(a[16]),
.I1(b[17]),
.I2(a[15]),
.I3(b[18]),
.I4(a[14]),
.I5(b[19]));

wire p_s0_o31_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v5 (
.O6(p_s0_o31_5),
.O5(),
.I0(a[16]),
.I1(b[17]),
.I2(a[15]),
.I3(b[18]),
.I4(a[14]),
.I5(b[19]));

wire p_s0_o30_16;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v6 (
.O6(p_s0_o30_16),
.O5(),
.I0(a[13]),
.I1(b[20]),
.I2(a[12]),
.I3(b[21]),
.I4(a[11]),
.I5(b[22]));

wire p_s0_o31_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v6 (
.O6(p_s0_o31_6),
.O5(),
.I0(a[13]),
.I1(b[20]),
.I2(a[12]),
.I3(b[21]),
.I4(a[11]),
.I5(b[22]));

wire p_s0_o30_17;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v7 (
.O6(p_s0_o30_17),
.O5(),
.I0(a[10]),
.I1(b[23]),
.I2(a[9]),
.I3(b[24]),
.I4(a[8]),
.I5(b[25]));

wire p_s0_o31_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v7 (
.O6(p_s0_o31_7),
.O5(),
.I0(a[10]),
.I1(b[23]),
.I2(a[9]),
.I3(b[24]),
.I4(a[8]),
.I5(b[25]));

wire p_s0_o30_18;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o30_t24_z0_v8 (
.O6(p_s0_o30_18),
.O5(),
.I0(a[7]),
.I1(b[26]),
.I2(a[6]),
.I3(b[27]),
.I4(a[5]),
.I5(b[28]));

wire p_s0_o31_8;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o30_t24_z1_v8 (
.O6(p_s0_o31_8),
.O5(),
.I0(a[7]),
.I1(b[26]),
.I2(a[6]),
.I3(b[27]),
.I4(a[5]),
.I5(b[28]));

/////////STEP0----ORDER31////////////

wire p_s0_o31_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v0 (
.O6(p_s0_o31_9),
.O5(),
.I0(a[31]),
.I1(b[3]),
.I2(a[30]),
.I3(b[4]),
.I4(a[29]),
.I5(b[5]));

wire p_s0_o32_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v0 (
.O6(p_s0_o32_0),
.O5(),
.I0(a[31]),
.I1(b[3]),
.I2(a[30]),
.I3(b[4]),
.I4(a[29]),
.I5(b[5]));

wire p_s0_o31_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v1 (
.O6(p_s0_o31_10),
.O5(),
.I0(a[28]),
.I1(b[6]),
.I2(a[27]),
.I3(b[7]),
.I4(a[26]),
.I5(b[8]));

wire p_s0_o32_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v1 (
.O6(p_s0_o32_1),
.O5(),
.I0(a[28]),
.I1(b[6]),
.I2(a[27]),
.I3(b[7]),
.I4(a[26]),
.I5(b[8]));

wire p_s0_o31_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v2 (
.O6(p_s0_o31_11),
.O5(),
.I0(a[25]),
.I1(b[9]),
.I2(a[24]),
.I3(b[10]),
.I4(a[23]),
.I5(b[11]));

wire p_s0_o32_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v2 (
.O6(p_s0_o32_2),
.O5(),
.I0(a[25]),
.I1(b[9]),
.I2(a[24]),
.I3(b[10]),
.I4(a[23]),
.I5(b[11]));

wire p_s0_o31_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v3 (
.O6(p_s0_o31_12),
.O5(),
.I0(a[22]),
.I1(b[12]),
.I2(a[21]),
.I3(b[13]),
.I4(a[20]),
.I5(b[14]));

wire p_s0_o32_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v3 (
.O6(p_s0_o32_3),
.O5(),
.I0(a[22]),
.I1(b[12]),
.I2(a[21]),
.I3(b[13]),
.I4(a[20]),
.I5(b[14]));

wire p_s0_o31_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v4 (
.O6(p_s0_o31_13),
.O5(),
.I0(a[19]),
.I1(b[15]),
.I2(a[18]),
.I3(b[16]),
.I4(a[17]),
.I5(b[17]));

wire p_s0_o32_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v4 (
.O6(p_s0_o32_4),
.O5(),
.I0(a[19]),
.I1(b[15]),
.I2(a[18]),
.I3(b[16]),
.I4(a[17]),
.I5(b[17]));

wire p_s0_o31_14;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v5 (
.O6(p_s0_o31_14),
.O5(),
.I0(a[16]),
.I1(b[18]),
.I2(a[15]),
.I3(b[19]),
.I4(a[14]),
.I5(b[20]));

wire p_s0_o32_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v5 (
.O6(p_s0_o32_5),
.O5(),
.I0(a[16]),
.I1(b[18]),
.I2(a[15]),
.I3(b[19]),
.I4(a[14]),
.I5(b[20]));

wire p_s0_o31_15;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v6 (
.O6(p_s0_o31_15),
.O5(),
.I0(a[13]),
.I1(b[21]),
.I2(a[12]),
.I3(b[22]),
.I4(a[11]),
.I5(b[23]));

wire p_s0_o32_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v6 (
.O6(p_s0_o32_6),
.O5(),
.I0(a[13]),
.I1(b[21]),
.I2(a[12]),
.I3(b[22]),
.I4(a[11]),
.I5(b[23]));

wire p_s0_o31_16;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v7 (
.O6(p_s0_o31_16),
.O5(),
.I0(a[10]),
.I1(b[24]),
.I2(a[9]),
.I3(b[25]),
.I4(a[8]),
.I5(b[26]));

wire p_s0_o32_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v7 (
.O6(p_s0_o32_7),
.O5(),
.I0(a[10]),
.I1(b[24]),
.I2(a[9]),
.I3(b[25]),
.I4(a[8]),
.I5(b[26]));

wire p_s0_o31_17;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o31_t25_z0_v8 (
.O6(p_s0_o31_17),
.O5(),
.I0(a[7]),
.I1(b[27]),
.I2(a[6]),
.I3(b[28]),
.I4(a[5]),
.I5(b[29]));

wire p_s0_o32_8;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o31_t25_z1_v8 (
.O6(p_s0_o32_8),
.O5(),
.I0(a[7]),
.I1(b[27]),
.I2(a[6]),
.I3(b[28]),
.I4(a[5]),
.I5(b[29]));

/////////STEP0----ORDER32////////////

wire p_s0_o32_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o32_t26_z0_v0 (
.O6(p_s0_o32_9),
.O5(),
.I0(a[31]),
.I1(b[4]),
.I2(a[30]),
.I3(b[5]),
.I4(a[29]),
.I5(b[6]));

wire p_s0_o33_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o32_t26_z1_v0 (
.O6(p_s0_o33_0),
.O5(),
.I0(a[31]),
.I1(b[4]),
.I2(a[30]),
.I3(b[5]),
.I4(a[29]),
.I5(b[6]));

wire p_s0_o32_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o32_t26_z0_v1 (
.O6(p_s0_o32_10),
.O5(),
.I0(a[28]),
.I1(b[7]),
.I2(a[27]),
.I3(b[8]),
.I4(a[26]),
.I5(b[9]));

wire p_s0_o33_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o32_t26_z1_v1 (
.O6(p_s0_o33_1),
.O5(),
.I0(a[28]),
.I1(b[7]),
.I2(a[27]),
.I3(b[8]),
.I4(a[26]),
.I5(b[9]));

wire p_s0_o32_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o32_t26_z0_v2 (
.O6(p_s0_o32_11),
.O5(),
.I0(a[25]),
.I1(b[10]),
.I2(a[24]),
.I3(b[11]),
.I4(a[23]),
.I5(b[12]));

wire p_s0_o33_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o32_t26_z1_v2 (
.O6(p_s0_o33_2),
.O5(),
.I0(a[25]),
.I1(b[10]),
.I2(a[24]),
.I3(b[11]),
.I4(a[23]),
.I5(b[12]));

wire p_s0_o32_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o32_t26_z0_v3 (
.O6(p_s0_o32_12),
.O5(),
.I0(a[22]),
.I1(b[13]),
.I2(a[21]),
.I3(b[14]),
.I4(a[20]),
.I5(b[15]));

wire p_s0_o33_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o32_t26_z1_v3 (
.O6(p_s0_o33_3),
.O5(),
.I0(a[22]),
.I1(b[13]),
.I2(a[21]),
.I3(b[14]),
.I4(a[20]),
.I5(b[15]));

wire p_s0_o32_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o32_t26_z0_v4 (
.O6(p_s0_o32_13),
.O5(),
.I0(a[19]),
.I1(b[16]),
.I2(a[18]),
.I3(b[17]),
.I4(a[17]),
.I5(b[18]));

wire p_s0_o33_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o32_t26_z1_v4 (
.O6(p_s0_o33_4),
.O5(),
.I0(a[19]),
.I1(b[16]),
.I2(a[18]),
.I3(b[17]),
.I4(a[17]),
.I5(b[18]));

wire p_s0_o32_14;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o32_t26_z0_v5 (
.O6(p_s0_o32_14),
.O5(),
.I0(a[16]),
.I1(b[19]),
.I2(a[15]),
.I3(b[20]),
.I4(a[14]),
.I5(b[21]));

wire p_s0_o33_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o32_t26_z1_v5 (
.O6(p_s0_o33_5),
.O5(),
.I0(a[16]),
.I1(b[19]),
.I2(a[15]),
.I3(b[20]),
.I4(a[14]),
.I5(b[21]));

wire p_s0_o32_15;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o32_t26_z0_v6 (
.O6(p_s0_o32_15),
.O5(),
.I0(a[13]),
.I1(b[22]),
.I2(a[12]),
.I3(b[23]),
.I4(a[11]),
.I5(b[24]));

wire p_s0_o33_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o32_t26_z1_v6 (
.O6(p_s0_o33_6),
.O5(),
.I0(a[13]),
.I1(b[22]),
.I2(a[12]),
.I3(b[23]),
.I4(a[11]),
.I5(b[24]));

wire p_s0_o32_16;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o32_t26_z0_v7 (
.O6(p_s0_o32_16),
.O5(),
.I0(a[10]),
.I1(b[25]),
.I2(a[9]),
.I3(b[26]),
.I4(a[8]),
.I5(b[27]));

wire p_s0_o33_7;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o32_t26_z1_v7 (
.O6(p_s0_o33_7),
.O5(),
.I0(a[10]),
.I1(b[25]),
.I2(a[9]),
.I3(b[26]),
.I4(a[8]),
.I5(b[27]));

/////////STEP0----ORDER33////////////

wire p_s0_o33_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o33_t27_z0_v0 (
.O6(p_s0_o33_8),
.O5(),
.I0(a[31]),
.I1(b[5]),
.I2(a[30]),
.I3(b[6]),
.I4(a[29]),
.I5(b[7]));

wire p_s0_o34_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o33_t27_z1_v0 (
.O6(p_s0_o34_0),
.O5(),
.I0(a[31]),
.I1(b[5]),
.I2(a[30]),
.I3(b[6]),
.I4(a[29]),
.I5(b[7]));

wire p_s0_o33_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o33_t27_z0_v1 (
.O6(p_s0_o33_9),
.O5(),
.I0(a[28]),
.I1(b[8]),
.I2(a[27]),
.I3(b[9]),
.I4(a[26]),
.I5(b[10]));

wire p_s0_o34_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o33_t27_z1_v1 (
.O6(p_s0_o34_1),
.O5(),
.I0(a[28]),
.I1(b[8]),
.I2(a[27]),
.I3(b[9]),
.I4(a[26]),
.I5(b[10]));

wire p_s0_o33_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o33_t27_z0_v2 (
.O6(p_s0_o33_10),
.O5(),
.I0(a[25]),
.I1(b[11]),
.I2(a[24]),
.I3(b[12]),
.I4(a[23]),
.I5(b[13]));

wire p_s0_o34_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o33_t27_z1_v2 (
.O6(p_s0_o34_2),
.O5(),
.I0(a[25]),
.I1(b[11]),
.I2(a[24]),
.I3(b[12]),
.I4(a[23]),
.I5(b[13]));

wire p_s0_o33_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o33_t27_z0_v3 (
.O6(p_s0_o33_11),
.O5(),
.I0(a[22]),
.I1(b[14]),
.I2(a[21]),
.I3(b[15]),
.I4(a[20]),
.I5(b[16]));

wire p_s0_o34_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o33_t27_z1_v3 (
.O6(p_s0_o34_3),
.O5(),
.I0(a[22]),
.I1(b[14]),
.I2(a[21]),
.I3(b[15]),
.I4(a[20]),
.I5(b[16]));

wire p_s0_o33_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o33_t27_z0_v4 (
.O6(p_s0_o33_12),
.O5(),
.I0(a[19]),
.I1(b[17]),
.I2(a[18]),
.I3(b[18]),
.I4(a[17]),
.I5(b[19]));

wire p_s0_o34_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o33_t27_z1_v4 (
.O6(p_s0_o34_4),
.O5(),
.I0(a[19]),
.I1(b[17]),
.I2(a[18]),
.I3(b[18]),
.I4(a[17]),
.I5(b[19]));

wire p_s0_o33_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o33_t27_z0_v5 (
.O6(p_s0_o33_13),
.O5(),
.I0(a[16]),
.I1(b[20]),
.I2(a[15]),
.I3(b[21]),
.I4(a[14]),
.I5(b[22]));

wire p_s0_o34_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o33_t27_z1_v5 (
.O6(p_s0_o34_5),
.O5(),
.I0(a[16]),
.I1(b[20]),
.I2(a[15]),
.I3(b[21]),
.I4(a[14]),
.I5(b[22]));

wire p_s0_o33_14;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o33_t27_z0_v6 (
.O6(p_s0_o33_14),
.O5(),
.I0(a[13]),
.I1(b[23]),
.I2(a[12]),
.I3(b[24]),
.I4(a[11]),
.I5(b[25]));

wire p_s0_o34_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o33_t27_z1_v6 (
.O6(p_s0_o34_6),
.O5(),
.I0(a[13]),
.I1(b[23]),
.I2(a[12]),
.I3(b[24]),
.I4(a[11]),
.I5(b[25]));

/////////STEP0----ORDER34////////////

wire p_s0_o34_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o34_t28_z0_v0 (
.O6(p_s0_o34_7),
.O5(),
.I0(a[31]),
.I1(b[6]),
.I2(a[30]),
.I3(b[7]),
.I4(a[29]),
.I5(b[8]));

wire p_s0_o35_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o34_t28_z1_v0 (
.O6(p_s0_o35_0),
.O5(),
.I0(a[31]),
.I1(b[6]),
.I2(a[30]),
.I3(b[7]),
.I4(a[29]),
.I5(b[8]));

wire p_s0_o34_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o34_t28_z0_v1 (
.O6(p_s0_o34_8),
.O5(),
.I0(a[28]),
.I1(b[9]),
.I2(a[27]),
.I3(b[10]),
.I4(a[26]),
.I5(b[11]));

wire p_s0_o35_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o34_t28_z1_v1 (
.O6(p_s0_o35_1),
.O5(),
.I0(a[28]),
.I1(b[9]),
.I2(a[27]),
.I3(b[10]),
.I4(a[26]),
.I5(b[11]));

wire p_s0_o34_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o34_t28_z0_v2 (
.O6(p_s0_o34_9),
.O5(),
.I0(a[25]),
.I1(b[12]),
.I2(a[24]),
.I3(b[13]),
.I4(a[23]),
.I5(b[14]));

wire p_s0_o35_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o34_t28_z1_v2 (
.O6(p_s0_o35_2),
.O5(),
.I0(a[25]),
.I1(b[12]),
.I2(a[24]),
.I3(b[13]),
.I4(a[23]),
.I5(b[14]));

wire p_s0_o34_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o34_t28_z0_v3 (
.O6(p_s0_o34_10),
.O5(),
.I0(a[22]),
.I1(b[15]),
.I2(a[21]),
.I3(b[16]),
.I4(a[20]),
.I5(b[17]));

wire p_s0_o35_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o34_t28_z1_v3 (
.O6(p_s0_o35_3),
.O5(),
.I0(a[22]),
.I1(b[15]),
.I2(a[21]),
.I3(b[16]),
.I4(a[20]),
.I5(b[17]));

wire p_s0_o34_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o34_t28_z0_v4 (
.O6(p_s0_o34_11),
.O5(),
.I0(a[19]),
.I1(b[18]),
.I2(a[18]),
.I3(b[19]),
.I4(a[17]),
.I5(b[20]));

wire p_s0_o35_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o34_t28_z1_v4 (
.O6(p_s0_o35_4),
.O5(),
.I0(a[19]),
.I1(b[18]),
.I2(a[18]),
.I3(b[19]),
.I4(a[17]),
.I5(b[20]));

wire p_s0_o34_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o34_t28_z0_v5 (
.O6(p_s0_o34_12),
.O5(),
.I0(a[16]),
.I1(b[21]),
.I2(a[15]),
.I3(b[22]),
.I4(a[14]),
.I5(b[23]));

wire p_s0_o35_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o34_t28_z1_v5 (
.O6(p_s0_o35_5),
.O5(),
.I0(a[16]),
.I1(b[21]),
.I2(a[15]),
.I3(b[22]),
.I4(a[14]),
.I5(b[23]));

wire p_s0_o34_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o34_t28_z0_v6 (
.O6(p_s0_o34_13),
.O5(),
.I0(a[13]),
.I1(b[24]),
.I2(a[12]),
.I3(b[25]),
.I4(a[11]),
.I5(b[26]));

wire p_s0_o35_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o34_t28_z1_v6 (
.O6(p_s0_o35_6),
.O5(),
.I0(a[13]),
.I1(b[24]),
.I2(a[12]),
.I3(b[25]),
.I4(a[11]),
.I5(b[26]));

/////////STEP0----ORDER35////////////

wire p_s0_o35_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o35_t29_z0_v0 (
.O6(p_s0_o35_7),
.O5(),
.I0(a[31]),
.I1(b[7]),
.I2(a[30]),
.I3(b[8]),
.I4(a[29]),
.I5(b[9]));

wire p_s0_o36_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o35_t29_z1_v0 (
.O6(p_s0_o36_0),
.O5(),
.I0(a[31]),
.I1(b[7]),
.I2(a[30]),
.I3(b[8]),
.I4(a[29]),
.I5(b[9]));

wire p_s0_o35_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o35_t29_z0_v1 (
.O6(p_s0_o35_8),
.O5(),
.I0(a[28]),
.I1(b[10]),
.I2(a[27]),
.I3(b[11]),
.I4(a[26]),
.I5(b[12]));

wire p_s0_o36_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o35_t29_z1_v1 (
.O6(p_s0_o36_1),
.O5(),
.I0(a[28]),
.I1(b[10]),
.I2(a[27]),
.I3(b[11]),
.I4(a[26]),
.I5(b[12]));

wire p_s0_o35_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o35_t29_z0_v2 (
.O6(p_s0_o35_9),
.O5(),
.I0(a[25]),
.I1(b[13]),
.I2(a[24]),
.I3(b[14]),
.I4(a[23]),
.I5(b[15]));

wire p_s0_o36_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o35_t29_z1_v2 (
.O6(p_s0_o36_2),
.O5(),
.I0(a[25]),
.I1(b[13]),
.I2(a[24]),
.I3(b[14]),
.I4(a[23]),
.I5(b[15]));

wire p_s0_o35_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o35_t29_z0_v3 (
.O6(p_s0_o35_10),
.O5(),
.I0(a[22]),
.I1(b[16]),
.I2(a[21]),
.I3(b[17]),
.I4(a[20]),
.I5(b[18]));

wire p_s0_o36_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o35_t29_z1_v3 (
.O6(p_s0_o36_3),
.O5(),
.I0(a[22]),
.I1(b[16]),
.I2(a[21]),
.I3(b[17]),
.I4(a[20]),
.I5(b[18]));

wire p_s0_o35_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o35_t29_z0_v4 (
.O6(p_s0_o35_11),
.O5(),
.I0(a[19]),
.I1(b[19]),
.I2(a[18]),
.I3(b[20]),
.I4(a[17]),
.I5(b[21]));

wire p_s0_o36_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o35_t29_z1_v4 (
.O6(p_s0_o36_4),
.O5(),
.I0(a[19]),
.I1(b[19]),
.I2(a[18]),
.I3(b[20]),
.I4(a[17]),
.I5(b[21]));

wire p_s0_o35_12;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o35_t29_z0_v5 (
.O6(p_s0_o35_12),
.O5(),
.I0(a[16]),
.I1(b[22]),
.I2(a[15]),
.I3(b[23]),
.I4(a[14]),
.I5(b[24]));

wire p_s0_o36_5;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o35_t29_z1_v5 (
.O6(p_s0_o36_5),
.O5(),
.I0(a[16]),
.I1(b[22]),
.I2(a[15]),
.I3(b[23]),
.I4(a[14]),
.I5(b[24]));

wire p_s0_o35_13;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o35_t29_z0_v6 (
.O6(p_s0_o35_13),
.O5(),
.I0(a[13]),
.I1(b[25]),
.I2(a[12]),
.I3(b[26]),
.I4(a[11]),
.I5(b[27]));

wire p_s0_o36_6;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o35_t29_z1_v6 (
.O6(p_s0_o36_6),
.O5(),
.I0(a[13]),
.I1(b[25]),
.I2(a[12]),
.I3(b[26]),
.I4(a[11]),
.I5(b[27]));

/////////STEP0----ORDER36////////////

wire p_s0_o36_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o36_t30_z0_v0 (
.O6(p_s0_o36_7),
.O5(),
.I0(a[31]),
.I1(b[8]),
.I2(a[30]),
.I3(b[9]),
.I4(a[29]),
.I5(b[10]));

wire p_s0_o37_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o36_t30_z1_v0 (
.O6(p_s0_o37_0),
.O5(),
.I0(a[31]),
.I1(b[8]),
.I2(a[30]),
.I3(b[9]),
.I4(a[29]),
.I5(b[10]));

wire p_s0_o36_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o36_t30_z0_v1 (
.O6(p_s0_o36_8),
.O5(),
.I0(a[28]),
.I1(b[11]),
.I2(a[27]),
.I3(b[12]),
.I4(a[26]),
.I5(b[13]));

wire p_s0_o37_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o36_t30_z1_v1 (
.O6(p_s0_o37_1),
.O5(),
.I0(a[28]),
.I1(b[11]),
.I2(a[27]),
.I3(b[12]),
.I4(a[26]),
.I5(b[13]));

wire p_s0_o36_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o36_t30_z0_v2 (
.O6(p_s0_o36_9),
.O5(),
.I0(a[25]),
.I1(b[14]),
.I2(a[24]),
.I3(b[15]),
.I4(a[23]),
.I5(b[16]));

wire p_s0_o37_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o36_t30_z1_v2 (
.O6(p_s0_o37_2),
.O5(),
.I0(a[25]),
.I1(b[14]),
.I2(a[24]),
.I3(b[15]),
.I4(a[23]),
.I5(b[16]));

wire p_s0_o36_10;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o36_t30_z0_v3 (
.O6(p_s0_o36_10),
.O5(),
.I0(a[22]),
.I1(b[17]),
.I2(a[21]),
.I3(b[18]),
.I4(a[20]),
.I5(b[19]));

wire p_s0_o37_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o36_t30_z1_v3 (
.O6(p_s0_o37_3),
.O5(),
.I0(a[22]),
.I1(b[17]),
.I2(a[21]),
.I3(b[18]),
.I4(a[20]),
.I5(b[19]));

wire p_s0_o36_11;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o36_t30_z0_v4 (
.O6(p_s0_o36_11),
.O5(),
.I0(a[19]),
.I1(b[20]),
.I2(a[18]),
.I3(b[21]),
.I4(a[17]),
.I5(b[22]));

wire p_s0_o37_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o36_t30_z1_v4 (
.O6(p_s0_o37_4),
.O5(),
.I0(a[19]),
.I1(b[20]),
.I2(a[18]),
.I3(b[21]),
.I4(a[17]),
.I5(b[22]));

/////////STEP0----ORDER37////////////

wire p_s0_o37_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o37_t31_z0_v0 (
.O6(p_s0_o37_5),
.O5(),
.I0(a[31]),
.I1(b[9]),
.I2(a[30]),
.I3(b[10]),
.I4(a[29]),
.I5(b[11]));

wire p_s0_o38_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o37_t31_z1_v0 (
.O6(p_s0_o38_0),
.O5(),
.I0(a[31]),
.I1(b[9]),
.I2(a[30]),
.I3(b[10]),
.I4(a[29]),
.I5(b[11]));

wire p_s0_o37_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o37_t31_z0_v1 (
.O6(p_s0_o37_6),
.O5(),
.I0(a[28]),
.I1(b[12]),
.I2(a[27]),
.I3(b[13]),
.I4(a[26]),
.I5(b[14]));

wire p_s0_o38_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o37_t31_z1_v1 (
.O6(p_s0_o38_1),
.O5(),
.I0(a[28]),
.I1(b[12]),
.I2(a[27]),
.I3(b[13]),
.I4(a[26]),
.I5(b[14]));

wire p_s0_o37_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o37_t31_z0_v2 (
.O6(p_s0_o37_7),
.O5(),
.I0(a[25]),
.I1(b[15]),
.I2(a[24]),
.I3(b[16]),
.I4(a[23]),
.I5(b[17]));

wire p_s0_o38_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o37_t31_z1_v2 (
.O6(p_s0_o38_2),
.O5(),
.I0(a[25]),
.I1(b[15]),
.I2(a[24]),
.I3(b[16]),
.I4(a[23]),
.I5(b[17]));

wire p_s0_o37_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o37_t31_z0_v3 (
.O6(p_s0_o37_8),
.O5(),
.I0(a[22]),
.I1(b[18]),
.I2(a[21]),
.I3(b[19]),
.I4(a[20]),
.I5(b[20]));

wire p_s0_o38_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o37_t31_z1_v3 (
.O6(p_s0_o38_3),
.O5(),
.I0(a[22]),
.I1(b[18]),
.I2(a[21]),
.I3(b[19]),
.I4(a[20]),
.I5(b[20]));

wire p_s0_o37_9;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o37_t31_z0_v4 (
.O6(p_s0_o37_9),
.O5(),
.I0(a[19]),
.I1(b[21]),
.I2(a[18]),
.I3(b[22]),
.I4(a[17]),
.I5(b[23]));

wire p_s0_o38_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o37_t31_z1_v4 (
.O6(p_s0_o38_4),
.O5(),
.I0(a[19]),
.I1(b[21]),
.I2(a[18]),
.I3(b[22]),
.I4(a[17]),
.I5(b[23]));

/////////STEP0----ORDER38////////////

wire p_s0_o38_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o38_t32_z0_v0 (
.O6(p_s0_o38_5),
.O5(),
.I0(a[31]),
.I1(b[10]),
.I2(a[30]),
.I3(b[11]),
.I4(a[29]),
.I5(b[12]));

wire p_s0_o39_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o38_t32_z1_v0 (
.O6(p_s0_o39_0),
.O5(),
.I0(a[31]),
.I1(b[10]),
.I2(a[30]),
.I3(b[11]),
.I4(a[29]),
.I5(b[12]));

wire p_s0_o38_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o38_t32_z0_v1 (
.O6(p_s0_o38_6),
.O5(),
.I0(a[28]),
.I1(b[13]),
.I2(a[27]),
.I3(b[14]),
.I4(a[26]),
.I5(b[15]));

wire p_s0_o39_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o38_t32_z1_v1 (
.O6(p_s0_o39_1),
.O5(),
.I0(a[28]),
.I1(b[13]),
.I2(a[27]),
.I3(b[14]),
.I4(a[26]),
.I5(b[15]));

wire p_s0_o38_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o38_t32_z0_v2 (
.O6(p_s0_o38_7),
.O5(),
.I0(a[25]),
.I1(b[16]),
.I2(a[24]),
.I3(b[17]),
.I4(a[23]),
.I5(b[18]));

wire p_s0_o39_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o38_t32_z1_v2 (
.O6(p_s0_o39_2),
.O5(),
.I0(a[25]),
.I1(b[16]),
.I2(a[24]),
.I3(b[17]),
.I4(a[23]),
.I5(b[18]));

wire p_s0_o38_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o38_t32_z0_v3 (
.O6(p_s0_o38_8),
.O5(),
.I0(a[22]),
.I1(b[19]),
.I2(a[21]),
.I3(b[20]),
.I4(a[20]),
.I5(b[21]));

wire p_s0_o39_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o38_t32_z1_v3 (
.O6(p_s0_o39_3),
.O5(),
.I0(a[22]),
.I1(b[19]),
.I2(a[21]),
.I3(b[20]),
.I4(a[20]),
.I5(b[21]));

/////////STEP0----ORDER39////////////

wire p_s0_o39_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o39_t33_z0_v0 (
.O6(p_s0_o39_4),
.O5(),
.I0(a[31]),
.I1(b[11]),
.I2(a[30]),
.I3(b[12]),
.I4(a[29]),
.I5(b[13]));

wire p_s0_o40_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o39_t33_z1_v0 (
.O6(p_s0_o40_0),
.O5(),
.I0(a[31]),
.I1(b[11]),
.I2(a[30]),
.I3(b[12]),
.I4(a[29]),
.I5(b[13]));

wire p_s0_o39_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o39_t33_z0_v1 (
.O6(p_s0_o39_5),
.O5(),
.I0(a[28]),
.I1(b[14]),
.I2(a[27]),
.I3(b[15]),
.I4(a[26]),
.I5(b[16]));

wire p_s0_o40_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o39_t33_z1_v1 (
.O6(p_s0_o40_1),
.O5(),
.I0(a[28]),
.I1(b[14]),
.I2(a[27]),
.I3(b[15]),
.I4(a[26]),
.I5(b[16]));

wire p_s0_o39_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o39_t33_z0_v2 (
.O6(p_s0_o39_6),
.O5(),
.I0(a[25]),
.I1(b[17]),
.I2(a[24]),
.I3(b[18]),
.I4(a[23]),
.I5(b[19]));

wire p_s0_o40_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o39_t33_z1_v2 (
.O6(p_s0_o40_2),
.O5(),
.I0(a[25]),
.I1(b[17]),
.I2(a[24]),
.I3(b[18]),
.I4(a[23]),
.I5(b[19]));

wire p_s0_o39_7;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o39_t33_z0_v3 (
.O6(p_s0_o39_7),
.O5(),
.I0(a[22]),
.I1(b[20]),
.I2(a[21]),
.I3(b[21]),
.I4(a[20]),
.I5(b[22]));

wire p_s0_o40_3;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o39_t33_z1_v3 (
.O6(p_s0_o40_3),
.O5(),
.I0(a[22]),
.I1(b[20]),
.I2(a[21]),
.I3(b[21]),
.I4(a[20]),
.I5(b[22]));

wire p_s0_o39_8;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o39_t33_z0_v4 (
.O6(p_s0_o39_8),
.O5(),
.I0(a[19]),
.I1(b[23]),
.I2(a[18]),
.I3(b[24]),
.I4(a[17]),
.I5(b[25]));

wire p_s0_o40_4;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o39_t33_z1_v4 (
.O6(p_s0_o40_4),
.O5(),
.I0(a[19]),
.I1(b[23]),
.I2(a[18]),
.I3(b[24]),
.I4(a[17]),
.I5(b[25]));

/////////STEP0----ORDER40////////////

wire p_s0_o40_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o40_t34_z0_v0 (
.O6(p_s0_o40_5),
.O5(),
.I0(a[31]),
.I1(b[12]),
.I2(a[30]),
.I3(b[13]),
.I4(a[29]),
.I5(b[14]));

wire p_s0_o41_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o40_t34_z1_v0 (
.O6(p_s0_o41_0),
.O5(),
.I0(a[31]),
.I1(b[12]),
.I2(a[30]),
.I3(b[13]),
.I4(a[29]),
.I5(b[14]));

wire p_s0_o40_6;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o40_t34_z0_v1 (
.O6(p_s0_o40_6),
.O5(),
.I0(a[28]),
.I1(b[15]),
.I2(a[27]),
.I3(b[16]),
.I4(a[26]),
.I5(b[17]));

wire p_s0_o41_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o40_t34_z1_v1 (
.O6(p_s0_o41_1),
.O5(),
.I0(a[28]),
.I1(b[15]),
.I2(a[27]),
.I3(b[16]),
.I4(a[26]),
.I5(b[17]));

/////////STEP0----ORDER41////////////

wire p_s0_o41_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o41_t35_z0_v0 (
.O6(p_s0_o41_2),
.O5(),
.I0(a[31]),
.I1(b[13]),
.I2(a[30]),
.I3(b[14]),
.I4(a[29]),
.I5(b[15]));

wire p_s0_o42_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o41_t35_z1_v0 (
.O6(p_s0_o42_0),
.O5(),
.I0(a[31]),
.I1(b[13]),
.I2(a[30]),
.I3(b[14]),
.I4(a[29]),
.I5(b[15]));

wire p_s0_o41_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o41_t35_z0_v1 (
.O6(p_s0_o41_3),
.O5(),
.I0(a[28]),
.I1(b[16]),
.I2(a[27]),
.I3(b[17]),
.I4(a[26]),
.I5(b[18]));

wire p_s0_o42_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o41_t35_z1_v1 (
.O6(p_s0_o42_1),
.O5(),
.I0(a[28]),
.I1(b[16]),
.I2(a[27]),
.I3(b[17]),
.I4(a[26]),
.I5(b[18]));

wire p_s0_o41_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o41_t35_z0_v2 (
.O6(p_s0_o41_4),
.O5(),
.I0(a[25]),
.I1(b[19]),
.I2(a[24]),
.I3(b[20]),
.I4(a[23]),
.I5(b[21]));

wire p_s0_o42_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o41_t35_z1_v2 (
.O6(p_s0_o42_2),
.O5(),
.I0(a[25]),
.I1(b[19]),
.I2(a[24]),
.I3(b[20]),
.I4(a[23]),
.I5(b[21]));

/////////STEP0----ORDER42////////////

wire p_s0_o42_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o42_t36_z0_v0 (
.O6(p_s0_o42_3),
.O5(),
.I0(a[31]),
.I1(b[14]),
.I2(a[30]),
.I3(b[15]),
.I4(a[29]),
.I5(b[16]));

wire p_s0_o43_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o42_t36_z1_v0 (
.O6(p_s0_o43_0),
.O5(),
.I0(a[31]),
.I1(b[14]),
.I2(a[30]),
.I3(b[15]),
.I4(a[29]),
.I5(b[16]));

wire p_s0_o42_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o42_t36_z0_v1 (
.O6(p_s0_o42_4),
.O5(),
.I0(a[28]),
.I1(b[17]),
.I2(a[27]),
.I3(b[18]),
.I4(a[26]),
.I5(b[19]));

wire p_s0_o43_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o42_t36_z1_v1 (
.O6(p_s0_o43_1),
.O5(),
.I0(a[28]),
.I1(b[17]),
.I2(a[27]),
.I3(b[18]),
.I4(a[26]),
.I5(b[19]));

wire p_s0_o42_5;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o42_t36_z0_v2 (
.O6(p_s0_o42_5),
.O5(),
.I0(a[25]),
.I1(b[20]),
.I2(a[24]),
.I3(b[21]),
.I4(a[23]),
.I5(b[22]));

wire p_s0_o43_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o42_t36_z1_v2 (
.O6(p_s0_o43_2),
.O5(),
.I0(a[25]),
.I1(b[20]),
.I2(a[24]),
.I3(b[21]),
.I4(a[23]),
.I5(b[22]));

/////////STEP0----ORDER43////////////

wire p_s0_o43_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o43_t37_z0_v0 (
.O6(p_s0_o43_3),
.O5(),
.I0(a[31]),
.I1(b[15]),
.I2(a[30]),
.I3(b[16]),
.I4(a[29]),
.I5(b[17]));

wire p_s0_o44_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o43_t37_z1_v0 (
.O6(p_s0_o44_0),
.O5(),
.I0(a[31]),
.I1(b[15]),
.I2(a[30]),
.I3(b[16]),
.I4(a[29]),
.I5(b[17]));

wire p_s0_o43_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o43_t37_z0_v1 (
.O6(p_s0_o43_4),
.O5(),
.I0(a[28]),
.I1(b[18]),
.I2(a[27]),
.I3(b[19]),
.I4(a[26]),
.I5(b[20]));

wire p_s0_o44_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o43_t37_z1_v1 (
.O6(p_s0_o44_1),
.O5(),
.I0(a[28]),
.I1(b[18]),
.I2(a[27]),
.I3(b[19]),
.I4(a[26]),
.I5(b[20]));

/////////STEP0----ORDER44////////////

wire p_s0_o44_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o44_t38_z0_v0 (
.O6(p_s0_o44_2),
.O5(),
.I0(a[31]),
.I1(b[16]),
.I2(a[30]),
.I3(b[17]),
.I4(a[29]),
.I5(b[18]));

wire p_s0_o45_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o44_t38_z1_v0 (
.O6(p_s0_o45_0),
.O5(),
.I0(a[31]),
.I1(b[16]),
.I2(a[30]),
.I3(b[17]),
.I4(a[29]),
.I5(b[18]));

wire p_s0_o44_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o44_t38_z0_v1 (
.O6(p_s0_o44_3),
.O5(),
.I0(a[28]),
.I1(b[19]),
.I2(a[27]),
.I3(b[20]),
.I4(a[26]),
.I5(b[21]));

wire p_s0_o45_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o44_t38_z1_v1 (
.O6(p_s0_o45_1),
.O5(),
.I0(a[28]),
.I1(b[19]),
.I2(a[27]),
.I3(b[20]),
.I4(a[26]),
.I5(b[21]));

wire p_s0_o44_4;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o44_t38_z0_v2 (
.O6(p_s0_o44_4),
.O5(),
.I0(a[25]),
.I1(b[22]),
.I2(a[24]),
.I3(b[23]),
.I4(a[23]),
.I5(b[24]));

wire p_s0_o45_2;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o44_t38_z1_v2 (
.O6(p_s0_o45_2),
.O5(),
.I0(a[25]),
.I1(b[22]),
.I2(a[24]),
.I3(b[23]),
.I4(a[23]),
.I5(b[24]));

/////////STEP0----ORDER45////////////

wire p_s0_o45_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o45_t39_z0_v0 (
.O6(p_s0_o45_3),
.O5(),
.I0(a[31]),
.I1(b[17]),
.I2(a[30]),
.I3(b[18]),
.I4(a[29]),
.I5(b[19]));

wire p_s0_o46_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o45_t39_z1_v0 (
.O6(p_s0_o46_0),
.O5(),
.I0(a[31]),
.I1(b[17]),
.I2(a[30]),
.I3(b[18]),
.I4(a[29]),
.I5(b[19]));

/////////STEP0----ORDER46////////////

wire p_s0_o46_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o46_t40_z0_v0 (
.O6(p_s0_o46_1),
.O5(),
.I0(a[31]),
.I1(b[18]),
.I2(a[30]),
.I3(b[19]),
.I4(a[29]),
.I5(b[20]));

wire p_s0_o47_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o46_t40_z1_v0 (
.O6(p_s0_o47_0),
.O5(),
.I0(a[31]),
.I1(b[18]),
.I2(a[30]),
.I3(b[19]),
.I4(a[29]),
.I5(b[20]));

wire p_s0_o46_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o46_t40_z0_v1 (
.O6(p_s0_o46_2),
.O5(),
.I0(a[28]),
.I1(b[21]),
.I2(a[27]),
.I3(b[22]),
.I4(a[26]),
.I5(b[23]));

wire p_s0_o47_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o46_t40_z1_v1 (
.O6(p_s0_o47_1),
.O5(),
.I0(a[28]),
.I1(b[21]),
.I2(a[27]),
.I3(b[22]),
.I4(a[26]),
.I5(b[23]));

/////////STEP0----ORDER47////////////

wire p_s0_o47_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o47_t41_z0_v0 (
.O6(p_s0_o47_2),
.O5(),
.I0(a[31]),
.I1(b[19]),
.I2(a[30]),
.I3(b[20]),
.I4(a[29]),
.I5(b[21]));

wire p_s0_o48_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o47_t41_z1_v0 (
.O6(p_s0_o48_0),
.O5(),
.I0(a[31]),
.I1(b[19]),
.I2(a[30]),
.I3(b[20]),
.I4(a[29]),
.I5(b[21]));

/////////STEP0----ORDER48////////////

wire p_s0_o48_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o48_t42_z0_v0 (
.O6(p_s0_o48_1),
.O5(),
.I0(a[31]),
.I1(b[20]),
.I2(a[30]),
.I3(b[21]),
.I4(a[29]),
.I5(b[22]));

wire p_s0_o49_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o48_t42_z1_v0 (
.O6(p_s0_o49_0),
.O5(),
.I0(a[31]),
.I1(b[20]),
.I2(a[30]),
.I3(b[21]),
.I4(a[29]),
.I5(b[22]));

wire p_s0_o48_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o48_t42_z0_v1 (
.O6(p_s0_o48_2),
.O5(),
.I0(a[28]),
.I1(b[23]),
.I2(a[27]),
.I3(b[24]),
.I4(a[26]),
.I5(b[25]));

wire p_s0_o49_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o48_t42_z1_v1 (
.O6(p_s0_o49_1),
.O5(),
.I0(a[28]),
.I1(b[23]),
.I2(a[27]),
.I3(b[24]),
.I4(a[26]),
.I5(b[25]));

/////////STEP0----ORDER49////////////

/////////STEP0----ORDER50////////////

wire p_s0_o50_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o50_t43_z0_v0 (
.O6(p_s0_o50_0),
.O5(),
.I0(a[31]),
.I1(b[22]),
.I2(a[30]),
.I3(b[23]),
.I4(a[29]),
.I5(b[24]));

wire p_s0_o51_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o50_t43_z1_v0 (
.O6(p_s0_o51_0),
.O5(),
.I0(a[31]),
.I1(b[22]),
.I2(a[30]),
.I3(b[23]),
.I4(a[29]),
.I5(b[24]));

/////////STEP0----ORDER51////////////

wire p_s0_o51_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o51_t44_z0_v0 (
.O6(p_s0_o51_1),
.O5(),
.I0(a[31]),
.I1(b[23]),
.I2(a[30]),
.I3(b[24]),
.I4(a[29]),
.I5(b[25]));

wire p_s0_o52_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o51_t44_z1_v0 (
.O6(p_s0_o52_0),
.O5(),
.I0(a[31]),
.I1(b[23]),
.I2(a[30]),
.I3(b[24]),
.I4(a[29]),
.I5(b[25]));

/////////STEP0----ORDER52////////////

/////////STEP0----ORDER53////////////

/////////STEP0----ORDER54////////////

wire p_s0_o54_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o54_t45_z0_v0 (
.O6(p_s0_o54_0),
.O5(),
.I0(a[31]),
.I1(b[26]),
.I2(a[30]),
.I3(b[27]),
.I4(a[29]),
.I5(b[28]));

wire p_s0_o55_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o54_t45_z1_v0 (
.O6(p_s0_o55_0),
.O5(),
.I0(a[31]),
.I1(b[26]),
.I2(a[30]),
.I3(b[27]),
.I4(a[29]),
.I5(b[28]));

/////////STEP0----ORDER55////////////

/////////STEP0----ORDER56////////////

/////////STEP0----ORDER57////////////

/////////STEP0----ORDER58////////////

/////////STEP0----ORDER59////////////

/////////STEP1----ORDER0////////////

/////////STEP1----ORDER1////////////

wire p_s1_o2_0;
wire p_s1_o1_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o1_t60_z0_v0 (
.O6(p_s1_o2_0),
.O5(p_s1_o1_0),
.I0(a[4]),
.I1(b[0]),
.I2(a[3]),
.I3(b[1]),
.I4(p_s0_o1_0),
.I5(1'b1));

/////////STEP1----ORDER2////////////

/////////STEP1----ORDER3////////////

wire p_s1_o4_0;
wire p_s1_o3_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o3_t61_z0_v0 (
.O6(p_s1_o4_0),
.O5(p_s1_o3_0),
.I0(a[3]),
.I1(b[3]),
.I2(a[2]),
.I3(b[4]),
.I4(p_s0_o3_0),
.I5(1'b1));

/////////STEP1----ORDER4////////////

wire p_s1_o5_0;
wire p_s1_o4_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o4_t62_z0_v0 (
.O6(p_s1_o5_0),
.O5(p_s1_o4_1),
.I0(a[4]),
.I1(b[3]),
.I2(a[3]),
.I3(b[4]),
.I4(p_s0_o4_0),
.I5(1'b1));

wire p_s1_o5_1;
wire p_s1_o4_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o4_t62_z0_v1 (
.O6(p_s1_o5_1),
.O5(p_s1_o4_2),
.I0(a[2]),
.I1(b[5]),
.I2(a[1]),
.I3(b[6]),
.I4(p_s0_o4_1),
.I5(1'b1));

/////////STEP1----ORDER5////////////

wire p_s1_o6_0;
wire p_s1_o5_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o5_t63_z0_v0 (
.O6(p_s1_o6_0),
.O5(p_s1_o5_2),
.I0(a[8]),
.I1(b[0]),
.I2(a[7]),
.I3(b[1]),
.I4(p_s0_o5_0),
.I5(1'b1));

/////////STEP1----ORDER6////////////

/////////STEP1----ORDER7////////////

wire p_s1_o8_0;
wire p_s1_o7_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o7_t64_z0_v0 (
.O6(p_s1_o8_0),
.O5(p_s1_o7_0),
.I0(a[4]),
.I1(b[6]),
.I2(a[3]),
.I3(b[7]),
.I4(p_s0_o7_0),
.I5(1'b1));

wire p_s1_o8_1;
wire p_s1_o7_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o7_t64_z0_v1 (
.O6(p_s1_o8_1),
.O5(p_s1_o7_1),
.I0(a[2]),
.I1(b[8]),
.I2(a[1]),
.I3(b[9]),
.I4(p_s0_o7_1),
.I5(1'b1));

/////////STEP1----ORDER8////////////

wire p_s1_o9_0;
wire p_s1_o8_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o8_t65_z0_v0 (
.O6(p_s1_o9_0),
.O5(p_s1_o8_2),
.I0(a[11]),
.I1(b[0]),
.I2(a[10]),
.I3(b[1]),
.I4(p_s0_o8_0),
.I5(1'b1));

wire p_s1_o9_1;
wire p_s1_o8_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o8_t65_z0_v1 (
.O6(p_s1_o9_1),
.O5(p_s1_o8_3),
.I0(a[9]),
.I1(b[2]),
.I2(a[8]),
.I3(b[3]),
.I4(p_s0_o8_1),
.I5(1'b1));

/////////STEP1----ORDER9////////////

wire p_s1_o10_0;
wire p_s1_o9_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o9_t66_z0_v0 (
.O6(p_s1_o10_0),
.O5(p_s1_o9_2),
.I0(a[9]),
.I1(b[3]),
.I2(a[8]),
.I3(b[4]),
.I4(p_s0_o9_0),
.I5(1'b1));

/////////STEP1----ORDER10////////////

wire p_s1_o11_0;
wire p_s1_o10_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o10_t67_z0_v0 (
.O6(p_s1_o11_0),
.O5(p_s1_o10_1),
.I0(a[7]),
.I1(b[6]),
.I2(a[6]),
.I3(b[7]),
.I4(p_s0_o10_0),
.I5(1'b1));

wire p_s1_o11_1;
wire p_s1_o10_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o10_t67_z0_v1 (
.O6(p_s1_o11_1),
.O5(p_s1_o10_2),
.I0(a[5]),
.I1(b[8]),
.I2(a[4]),
.I3(b[9]),
.I4(p_s0_o10_1),
.I5(1'b1));

wire p_s1_o11_2;
wire p_s1_o10_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o10_t67_z0_v2 (
.O6(p_s1_o11_2),
.O5(p_s1_o10_3),
.I0(a[3]),
.I1(b[10]),
.I2(a[2]),
.I3(b[11]),
.I4(p_s0_o10_2),
.I5(1'b1));

/////////STEP1----ORDER11////////////

wire p_s1_o12_0;
wire p_s1_o11_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o11_t68_z0_v0 (
.O6(p_s1_o12_0),
.O5(p_s1_o11_3),
.I0(a[9]),
.I1(b[5]),
.I2(a[8]),
.I3(b[6]),
.I4(p_s0_o11_0),
.I5(1'b1));

wire p_s1_o12_1;
wire p_s1_o11_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o11_t68_z0_v1 (
.O6(p_s1_o12_1),
.O5(p_s1_o11_4),
.I0(a[7]),
.I1(b[7]),
.I2(a[6]),
.I3(b[8]),
.I4(p_s0_o11_1),
.I5(1'b1));

wire p_s1_o12_2;
wire p_s1_o11_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o11_t68_z0_v2 (
.O6(p_s1_o12_2),
.O5(p_s1_o11_5),
.I0(a[5]),
.I1(b[9]),
.I2(a[4]),
.I3(b[10]),
.I4(p_s0_o11_2),
.I5(1'b1));

wire p_s1_o12_3;
wire p_s1_o11_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o11_t68_z0_v3 (
.O6(p_s1_o12_3),
.O5(p_s1_o11_6),
.I0(a[3]),
.I1(b[11]),
.I2(a[2]),
.I3(b[12]),
.I4(p_s0_o11_3),
.I5(1'b1));

/////////STEP1----ORDER12////////////

wire p_s1_o13_0;
wire p_s1_o12_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o12_t69_z0_v0 (
.O6(p_s1_o13_0),
.O5(p_s1_o12_4),
.I0(a[13]),
.I1(b[2]),
.I2(a[12]),
.I3(b[3]),
.I4(p_s0_o12_0),
.I5(1'b1));

wire p_s1_o13_1;
wire p_s1_o12_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o12_t69_z0_v1 (
.O6(p_s1_o13_1),
.O5(p_s1_o12_5),
.I0(a[11]),
.I1(b[4]),
.I2(a[10]),
.I3(b[5]),
.I4(p_s0_o12_1),
.I5(1'b1));

wire p_s1_o13_2;
wire p_s1_o12_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o12_t69_z0_v2 (
.O6(p_s1_o13_2),
.O5(p_s1_o12_6),
.I0(a[9]),
.I1(b[6]),
.I2(a[8]),
.I3(b[7]),
.I4(p_s0_o12_2),
.I5(1'b1));

/////////STEP1----ORDER13////////////

wire p_s1_o14_0;
wire p_s1_o13_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o13_t70_z0_v0 (
.O6(p_s1_o14_0),
.O5(p_s1_o13_3),
.I0(a[1]),
.I1(b[15]),
.I2(a[0]),
.I3(b[16]),
.I4(p_s0_o13_0),
.I5(1'b1));

wire p_s1_o14_1;
wire p_s1_o13_4;
LUT6_2 #(
.INIT(64'h177E7EE896696996)
) LUT6_2_inst_s1_o13_t124_z0_v0 (
.O6(p_s1_o14_1),
.O5(p_s1_o13_4),
.I0(p_s0_o13_1),
.I1(p_s0_o13_2),
.I2(p_s0_o13_3),
.I3(p_s0_o13_4),
.I4(p_s0_o13_5),
.I5(1'b1));

wire p_s1_o15_0;
LUT6_2 #(
.INIT(64'hE8808000E8808000)
) LUT6_2_inst_s1_o13_t124_z1_v0 (
.O6(p_s1_o15_0),
.O5(),
.I0(p_s0_o13_1),
.I1(p_s0_o13_2),
.I2(p_s0_o13_3),
.I3(p_s0_o13_4),
.I4(p_s0_o13_5),
.I5(1'b1));

/////////STEP1----ORDER14////////////

wire p_s1_o15_1;
wire p_s1_o14_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t71_z0_v0 (
.O6(p_s1_o15_1),
.O5(p_s1_o14_2),
.I0(a[11]),
.I1(b[6]),
.I2(a[10]),
.I3(b[7]),
.I4(p_s0_o14_0),
.I5(1'b1));

wire p_s1_o15_2;
wire p_s1_o14_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t71_z0_v1 (
.O6(p_s1_o15_2),
.O5(p_s1_o14_3),
.I0(a[9]),
.I1(b[8]),
.I2(a[8]),
.I3(b[9]),
.I4(p_s0_o14_1),
.I5(1'b1));

wire p_s1_o15_3;
wire p_s1_o14_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t71_z0_v2 (
.O6(p_s1_o15_3),
.O5(p_s1_o14_4),
.I0(a[7]),
.I1(b[10]),
.I2(a[6]),
.I3(b[11]),
.I4(p_s0_o14_2),
.I5(1'b1));

wire p_s1_o15_4;
wire p_s1_o14_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t71_z0_v3 (
.O6(p_s1_o15_4),
.O5(p_s1_o14_5),
.I0(a[5]),
.I1(b[12]),
.I2(a[4]),
.I3(b[13]),
.I4(p_s0_o14_3),
.I5(1'b1));

wire p_s1_o15_5;
wire p_s1_o14_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t71_z0_v4 (
.O6(p_s1_o15_5),
.O5(p_s1_o14_6),
.I0(a[3]),
.I1(b[14]),
.I2(a[2]),
.I3(b[15]),
.I4(p_s0_o14_4),
.I5(1'b1));

wire p_s1_o15_6;
wire p_s1_o14_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t71_z0_v5 (
.O6(p_s1_o15_6),
.O5(p_s1_o14_7),
.I0(a[1]),
.I1(b[16]),
.I2(a[0]),
.I3(b[17]),
.I4(p_s0_o14_5),
.I5(1'b1));

/////////STEP1----ORDER15////////////

wire p_s1_o16_0;
wire p_s1_o15_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o15_t72_z0_v0 (
.O6(p_s1_o16_0),
.O5(p_s1_o15_7),
.I0(a[9]),
.I1(b[9]),
.I2(a[8]),
.I3(b[10]),
.I4(p_s0_o15_0),
.I5(1'b1));

wire p_s1_o16_1;
wire p_s1_o15_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o15_t72_z0_v1 (
.O6(p_s1_o16_1),
.O5(p_s1_o15_8),
.I0(a[7]),
.I1(b[11]),
.I2(a[6]),
.I3(b[12]),
.I4(p_s0_o15_1),
.I5(1'b1));

wire p_s1_o16_2;
wire p_s1_o15_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o15_t72_z0_v2 (
.O6(p_s1_o16_2),
.O5(p_s1_o15_9),
.I0(a[5]),
.I1(b[13]),
.I2(a[4]),
.I3(b[14]),
.I4(p_s0_o15_2),
.I5(1'b1));

wire p_s1_o16_3;
wire p_s1_o15_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o15_t72_z0_v3 (
.O6(p_s1_o16_3),
.O5(p_s1_o15_10),
.I0(a[3]),
.I1(b[15]),
.I2(a[2]),
.I3(b[16]),
.I4(p_s0_o15_3),
.I5(1'b1));

wire p_s1_o16_4;
wire p_s1_o15_11;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o15_t72_z0_v4 (
.O6(p_s1_o16_4),
.O5(p_s1_o15_11),
.I0(a[1]),
.I1(b[17]),
.I2(a[0]),
.I3(b[18]),
.I4(p_s0_o15_4),
.I5(1'b1));

/////////STEP1----ORDER16////////////

wire p_s1_o17_0;
wire p_s1_o16_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o16_t73_z0_v0 (
.O6(p_s1_o17_0),
.O5(p_s1_o16_5),
.I0(a[10]),
.I1(b[9]),
.I2(a[9]),
.I3(b[10]),
.I4(p_s0_o16_0),
.I5(1'b1));

wire p_s1_o17_1;
wire p_s1_o16_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o16_t73_z0_v1 (
.O6(p_s1_o17_1),
.O5(p_s1_o16_6),
.I0(a[8]),
.I1(b[11]),
.I2(a[7]),
.I3(b[12]),
.I4(p_s0_o16_1),
.I5(1'b1));

wire p_s1_o17_2;
wire p_s1_o16_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o16_t73_z0_v2 (
.O6(p_s1_o17_2),
.O5(p_s1_o16_7),
.I0(a[6]),
.I1(b[13]),
.I2(a[5]),
.I3(b[14]),
.I4(p_s0_o16_2),
.I5(1'b1));

wire p_s1_o17_3;
wire p_s1_o16_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o16_t73_z0_v3 (
.O6(p_s1_o17_3),
.O5(p_s1_o16_8),
.I0(a[4]),
.I1(b[15]),
.I2(a[3]),
.I3(b[16]),
.I4(p_s0_o16_3),
.I5(1'b1));

wire p_s1_o17_4;
wire p_s1_o16_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o16_t73_z0_v4 (
.O6(p_s1_o17_4),
.O5(p_s1_o16_9),
.I0(a[2]),
.I1(b[17]),
.I2(a[1]),
.I3(b[18]),
.I4(p_s0_o16_4),
.I5(1'b1));

/////////STEP1----ORDER17////////////

wire p_s1_o18_0;
wire p_s1_o17_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o17_t74_z0_v0 (
.O6(p_s1_o18_0),
.O5(p_s1_o17_5),
.I0(a[11]),
.I1(b[9]),
.I2(a[10]),
.I3(b[10]),
.I4(p_s0_o17_0),
.I5(1'b1));

wire p_s1_o18_1;
wire p_s1_o17_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o17_t74_z0_v1 (
.O6(p_s1_o18_1),
.O5(p_s1_o17_6),
.I0(a[9]),
.I1(b[11]),
.I2(a[8]),
.I3(b[12]),
.I4(p_s0_o17_1),
.I5(1'b1));

wire p_s1_o18_2;
wire p_s1_o17_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o17_t74_z0_v2 (
.O6(p_s1_o18_2),
.O5(p_s1_o17_7),
.I0(a[7]),
.I1(b[13]),
.I2(a[6]),
.I3(b[14]),
.I4(p_s0_o17_2),
.I5(1'b1));

wire p_s1_o18_3;
wire p_s1_o17_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o17_t74_z0_v3 (
.O6(p_s1_o18_3),
.O5(p_s1_o17_8),
.I0(a[5]),
.I1(b[15]),
.I2(a[4]),
.I3(b[16]),
.I4(p_s0_o17_3),
.I5(1'b1));

wire p_s1_o18_4;
wire p_s1_o17_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o17_t74_z0_v4 (
.O6(p_s1_o18_4),
.O5(p_s1_o17_9),
.I0(a[3]),
.I1(b[17]),
.I2(a[2]),
.I3(b[18]),
.I4(p_s0_o17_4),
.I5(1'b1));

wire p_s1_o18_5;
wire p_s1_o17_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o17_t74_z0_v5 (
.O6(p_s1_o18_5),
.O5(p_s1_o17_10),
.I0(a[1]),
.I1(b[19]),
.I2(a[0]),
.I3(b[20]),
.I4(p_s0_o17_5),
.I5(1'b1));

/////////STEP1----ORDER18////////////

wire p_s1_o19_0;
wire p_s1_o18_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o18_t75_z0_v0 (
.O6(p_s1_o19_0),
.O5(p_s1_o18_6),
.I0(a[9]),
.I1(b[12]),
.I2(a[8]),
.I3(b[13]),
.I4(p_s0_o18_0),
.I5(1'b1));

wire p_s1_o19_1;
wire p_s1_o18_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o18_t75_z0_v1 (
.O6(p_s1_o19_1),
.O5(p_s1_o18_7),
.I0(a[7]),
.I1(b[14]),
.I2(a[6]),
.I3(b[15]),
.I4(p_s0_o18_1),
.I5(1'b1));

wire p_s1_o19_2;
wire p_s1_o18_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o18_t75_z0_v2 (
.O6(p_s1_o19_2),
.O5(p_s1_o18_8),
.I0(a[5]),
.I1(b[16]),
.I2(a[4]),
.I3(b[17]),
.I4(p_s0_o18_2),
.I5(1'b1));

wire p_s1_o19_3;
wire p_s1_o18_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o18_t75_z0_v3 (
.O6(p_s1_o19_3),
.O5(p_s1_o18_9),
.I0(a[3]),
.I1(b[18]),
.I2(a[2]),
.I3(b[19]),
.I4(p_s0_o18_3),
.I5(1'b1));

wire p_s1_o19_4;
wire p_s1_o18_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o18_t75_z0_v4 (
.O6(p_s1_o19_4),
.O5(p_s1_o18_10),
.I0(a[1]),
.I1(b[20]),
.I2(a[0]),
.I3(b[21]),
.I4(p_s0_o18_4),
.I5(1'b1));

/////////STEP1----ORDER19////////////

wire p_s1_o20_0;
wire p_s1_o19_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t76_z0_v0 (
.O6(p_s1_o20_0),
.O5(p_s1_o19_5),
.I0(a[13]),
.I1(b[9]),
.I2(a[12]),
.I3(b[10]),
.I4(p_s0_o19_0),
.I5(1'b1));

wire p_s1_o20_1;
wire p_s1_o19_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t76_z0_v1 (
.O6(p_s1_o20_1),
.O5(p_s1_o19_6),
.I0(a[11]),
.I1(b[11]),
.I2(a[10]),
.I3(b[12]),
.I4(p_s0_o19_1),
.I5(1'b1));

wire p_s1_o20_2;
wire p_s1_o19_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t76_z0_v2 (
.O6(p_s1_o20_2),
.O5(p_s1_o19_7),
.I0(a[9]),
.I1(b[13]),
.I2(a[8]),
.I3(b[14]),
.I4(p_s0_o19_2),
.I5(1'b1));

wire p_s1_o20_3;
wire p_s1_o19_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t76_z0_v3 (
.O6(p_s1_o20_3),
.O5(p_s1_o19_8),
.I0(a[7]),
.I1(b[15]),
.I2(a[6]),
.I3(b[16]),
.I4(p_s0_o19_3),
.I5(1'b1));

wire p_s1_o20_4;
wire p_s1_o19_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t76_z0_v4 (
.O6(p_s1_o20_4),
.O5(p_s1_o19_9),
.I0(a[5]),
.I1(b[17]),
.I2(a[4]),
.I3(b[18]),
.I4(p_s0_o19_4),
.I5(1'b1));

wire p_s1_o20_5;
wire p_s1_o19_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t76_z0_v5 (
.O6(p_s1_o20_5),
.O5(p_s1_o19_10),
.I0(a[3]),
.I1(b[19]),
.I2(a[2]),
.I3(b[20]),
.I4(p_s0_o19_5),
.I5(1'b1));

wire p_s1_o20_6;
wire p_s1_o19_11;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t76_z0_v6 (
.O6(p_s1_o20_6),
.O5(p_s1_o19_11),
.I0(a[1]),
.I1(b[21]),
.I2(a[0]),
.I3(b[22]),
.I4(p_s0_o19_6),
.I5(1'b1));

/////////STEP1----ORDER20////////////

wire p_s1_o21_0;
wire p_s1_o20_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o20_t77_z0_v0 (
.O6(p_s1_o21_0),
.O5(p_s1_o20_7),
.I0(a[5]),
.I1(b[18]),
.I2(a[4]),
.I3(b[19]),
.I4(p_s0_o20_0),
.I5(1'b1));

wire p_s1_o21_1;
wire p_s1_o20_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o20_t77_z0_v1 (
.O6(p_s1_o21_1),
.O5(p_s1_o20_8),
.I0(a[3]),
.I1(b[20]),
.I2(a[2]),
.I3(b[21]),
.I4(p_s0_o20_1),
.I5(1'b1));

wire p_s1_o21_2;
wire p_s1_o20_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o20_t77_z0_v2 (
.O6(p_s1_o21_2),
.O5(p_s1_o20_9),
.I0(a[1]),
.I1(b[22]),
.I2(a[0]),
.I3(b[23]),
.I4(p_s0_o20_2),
.I5(1'b1));

wire p_s1_o21_3;
wire p_s1_o20_10;
LUT6_2 #(
.INIT(64'h81177EE869966996)
) LUT6_2_inst_s1_o20_t125_z0_v0 (
.O6(p_s1_o21_3),
.O5(p_s1_o20_10),
.I0(p_s0_o20_3),
.I1(p_s0_o20_4),
.I2(p_s0_o20_5),
.I3(p_s0_o20_6),
.I4(p_s0_o21_0),
.I5(1'b1));

wire p_s1_o22_0;
LUT6_2 #(
.INIT(64'hFEE88000FEE88000)
) LUT6_2_inst_s1_o20_t125_z1_v0 (
.O6(p_s1_o22_0),
.O5(),
.I0(p_s0_o20_3),
.I1(p_s0_o20_4),
.I2(p_s0_o20_5),
.I3(p_s0_o20_6),
.I4(p_s0_o21_0),
.I5(1'b1));

/////////STEP1----ORDER21////////////

wire p_s1_o22_1;
wire p_s1_o21_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o21_t78_z0_v0 (
.O6(p_s1_o22_1),
.O5(p_s1_o21_4),
.I0(a[15]),
.I1(b[9]),
.I2(a[14]),
.I3(b[10]),
.I4(p_s0_o21_1),
.I5(1'b1));

wire p_s1_o22_2;
wire p_s1_o21_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o21_t78_z0_v1 (
.O6(p_s1_o22_2),
.O5(p_s1_o21_5),
.I0(a[13]),
.I1(b[11]),
.I2(a[12]),
.I3(b[12]),
.I4(p_s0_o21_2),
.I5(1'b1));

wire p_s1_o22_3;
wire p_s1_o21_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o21_t78_z0_v2 (
.O6(p_s1_o22_3),
.O5(p_s1_o21_6),
.I0(a[11]),
.I1(b[13]),
.I2(a[10]),
.I3(b[14]),
.I4(p_s0_o21_3),
.I5(1'b1));

wire p_s1_o22_4;
wire p_s1_o21_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o21_t78_z0_v3 (
.O6(p_s1_o22_4),
.O5(p_s1_o21_7),
.I0(a[9]),
.I1(b[15]),
.I2(a[8]),
.I3(b[16]),
.I4(p_s0_o21_4),
.I5(1'b1));

wire p_s1_o22_5;
wire p_s1_o21_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o21_t78_z0_v4 (
.O6(p_s1_o22_5),
.O5(p_s1_o21_8),
.I0(a[7]),
.I1(b[17]),
.I2(a[6]),
.I3(b[18]),
.I4(p_s0_o21_5),
.I5(1'b1));

wire p_s1_o22_6;
wire p_s1_o21_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o21_t78_z0_v5 (
.O6(p_s1_o22_6),
.O5(p_s1_o21_9),
.I0(a[5]),
.I1(b[19]),
.I2(a[4]),
.I3(b[20]),
.I4(p_s0_o21_6),
.I5(1'b1));

wire p_s1_o22_7;
wire p_s1_o21_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o21_t78_z0_v6 (
.O6(p_s1_o22_7),
.O5(p_s1_o21_10),
.I0(a[3]),
.I1(b[21]),
.I2(a[2]),
.I3(b[22]),
.I4(p_s0_o21_7),
.I5(1'b1));

wire p_s1_o22_8;
wire p_s1_o21_11;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o21_t78_z0_v7 (
.O6(p_s1_o22_8),
.O5(p_s1_o21_11),
.I0(a[1]),
.I1(b[23]),
.I2(a[0]),
.I3(b[24]),
.I4(p_s0_o21_8),
.I5(1'b1));

/////////STEP1----ORDER22////////////

wire p_s1_o23_0;
wire p_s1_o22_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o22_t79_z0_v0 (
.O6(p_s1_o23_0),
.O5(p_s1_o22_9),
.I0(a[1]),
.I1(b[24]),
.I2(a[0]),
.I3(b[25]),
.I4(p_s0_o22_0),
.I5(1'b1));

wire p_s1_o22_10;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o22_t110_z0_v0 (
.O6(p_s1_o22_10),
.O5(),
.I0(p_s0_o22_1),
.I1(p_s0_o22_2),
.I2(p_s0_o22_3),
.I3(p_s0_o22_4),
.I4(p_s0_o22_5),
.I5(p_s0_o23_0));

wire p_s1_o23_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o22_t110_z1_v0 (
.O6(p_s1_o23_1),
.O5(),
.I0(p_s0_o22_1),
.I1(p_s0_o22_2),
.I2(p_s0_o22_3),
.I3(p_s0_o22_4),
.I4(p_s0_o22_5),
.I5(p_s0_o23_0));

wire p_s1_o24_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o22_t110_z2_v0 (
.O6(p_s1_o24_0),
.O5(),
.I0(p_s0_o22_1),
.I1(p_s0_o22_2),
.I2(p_s0_o22_3),
.I3(p_s0_o22_4),
.I4(p_s0_o22_5),
.I5(p_s0_o23_0));

wire p_s1_o22_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o22_t110_z0_v1 (
.O6(p_s1_o22_11),
.O5(),
.I0(p_s0_o22_6),
.I1(p_s0_o22_7),
.I2(p_s0_o22_8),
.I3(p_s0_o22_9),
.I4(p_s0_o22_10),
.I5(p_s0_o23_1));

wire p_s1_o23_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o22_t110_z1_v1 (
.O6(p_s1_o23_2),
.O5(),
.I0(p_s0_o22_6),
.I1(p_s0_o22_7),
.I2(p_s0_o22_8),
.I3(p_s0_o22_9),
.I4(p_s0_o22_10),
.I5(p_s0_o23_1));

wire p_s1_o24_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o22_t110_z2_v1 (
.O6(p_s1_o24_1),
.O5(),
.I0(p_s0_o22_6),
.I1(p_s0_o22_7),
.I2(p_s0_o22_8),
.I3(p_s0_o22_9),
.I4(p_s0_o22_10),
.I5(p_s0_o23_1));

/////////STEP1----ORDER23////////////

wire p_s1_o24_2;
wire p_s1_o23_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o23_t80_z0_v0 (
.O6(p_s1_o24_2),
.O5(p_s1_o23_3),
.I0(a[11]),
.I1(b[15]),
.I2(a[10]),
.I3(b[16]),
.I4(p_s0_o23_2),
.I5(1'b1));

wire p_s1_o24_3;
wire p_s1_o23_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o23_t80_z0_v1 (
.O6(p_s1_o24_3),
.O5(p_s1_o23_4),
.I0(a[9]),
.I1(b[17]),
.I2(a[8]),
.I3(b[18]),
.I4(p_s0_o23_3),
.I5(1'b1));

wire p_s1_o24_4;
wire p_s1_o23_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o23_t80_z0_v2 (
.O6(p_s1_o24_4),
.O5(p_s1_o23_5),
.I0(a[7]),
.I1(b[19]),
.I2(a[6]),
.I3(b[20]),
.I4(p_s0_o23_4),
.I5(1'b1));

wire p_s1_o24_5;
wire p_s1_o23_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o23_t80_z0_v3 (
.O6(p_s1_o24_5),
.O5(p_s1_o23_6),
.I0(a[5]),
.I1(b[21]),
.I2(a[4]),
.I3(b[22]),
.I4(p_s0_o23_5),
.I5(1'b1));

wire p_s1_o24_6;
wire p_s1_o23_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o23_t80_z0_v4 (
.O6(p_s1_o24_6),
.O5(p_s1_o23_7),
.I0(a[3]),
.I1(b[23]),
.I2(a[2]),
.I3(b[24]),
.I4(p_s0_o23_6),
.I5(1'b1));

wire p_s1_o24_7;
wire p_s1_o23_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o23_t80_z0_v5 (
.O6(p_s1_o24_7),
.O5(p_s1_o23_8),
.I0(a[1]),
.I1(b[25]),
.I2(a[0]),
.I3(b[26]),
.I4(p_s0_o23_7),
.I5(1'b1));

wire p_s1_o23_9;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o23_t111_z0_v0 (
.O6(p_s1_o23_9),
.O5(),
.I0(p_s0_o23_8),
.I1(p_s0_o23_9),
.I2(p_s0_o23_10),
.I3(p_s0_o23_11),
.I4(p_s0_o23_12),
.I5(p_s0_o24_0));

wire p_s1_o24_8;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o23_t111_z1_v0 (
.O6(p_s1_o24_8),
.O5(),
.I0(p_s0_o23_8),
.I1(p_s0_o23_9),
.I2(p_s0_o23_10),
.I3(p_s0_o23_11),
.I4(p_s0_o23_12),
.I5(p_s0_o24_0));

wire p_s1_o25_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o23_t111_z2_v0 (
.O6(p_s1_o25_0),
.O5(),
.I0(p_s0_o23_8),
.I1(p_s0_o23_9),
.I2(p_s0_o23_10),
.I3(p_s0_o23_11),
.I4(p_s0_o23_12),
.I5(p_s0_o24_0));

/////////STEP1----ORDER24////////////

wire p_s1_o25_1;
wire p_s1_o24_9;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o24_t51_z0_v0 (
.O6(p_s1_o25_1),
.O5(p_s1_o24_9),
.I0(a[0]),
.I1(b[27]),
.I2(p_s0_o24_1),
.I3(p_s0_o24_2),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o24_10;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s1_o24_t108_z0_v0 (
.O6(p_s1_o24_10),
.O5(),
.I0(p_s0_o24_3),
.I1(p_s0_o24_4),
.I2(p_s0_o24_5),
.I3(p_s0_o24_6),
.I4(p_s0_o24_7),
.I5(p_s0_o24_8));

wire p_s1_o25_2;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s1_o24_t108_z1_v0 (
.O6(p_s1_o25_2),
.O5(),
.I0(p_s0_o24_3),
.I1(p_s0_o24_4),
.I2(p_s0_o24_5),
.I3(p_s0_o24_6),
.I4(p_s0_o24_7),
.I5(p_s0_o24_8));

wire p_s1_o26_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s1_o24_t108_z2_v0 (
.O6(p_s1_o26_0),
.O5(),
.I0(p_s0_o24_3),
.I1(p_s0_o24_4),
.I2(p_s0_o24_5),
.I3(p_s0_o24_6),
.I4(p_s0_o24_7),
.I5(p_s0_o24_8));

wire p_s1_o24_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o24_t112_z0_v0 (
.O6(p_s1_o24_11),
.O5(),
.I0(p_s0_o24_9),
.I1(p_s0_o24_10),
.I2(p_s0_o24_11),
.I3(p_s0_o24_12),
.I4(p_s0_o24_13),
.I5(p_s0_o25_0));

wire p_s1_o25_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o24_t112_z1_v0 (
.O6(p_s1_o25_3),
.O5(),
.I0(p_s0_o24_9),
.I1(p_s0_o24_10),
.I2(p_s0_o24_11),
.I3(p_s0_o24_12),
.I4(p_s0_o24_13),
.I5(p_s0_o25_0));

wire p_s1_o26_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o24_t112_z2_v0 (
.O6(p_s1_o26_1),
.O5(),
.I0(p_s0_o24_9),
.I1(p_s0_o24_10),
.I2(p_s0_o24_11),
.I3(p_s0_o24_12),
.I4(p_s0_o24_13),
.I5(p_s0_o25_0));

/////////STEP1----ORDER25////////////

wire p_s1_o26_2;
wire p_s1_o25_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v0 (
.O6(p_s1_o26_2),
.O5(p_s1_o25_4),
.I0(a[19]),
.I1(b[9]),
.I2(a[18]),
.I3(b[10]),
.I4(p_s0_o25_1),
.I5(1'b1));

wire p_s1_o26_3;
wire p_s1_o25_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v1 (
.O6(p_s1_o26_3),
.O5(p_s1_o25_5),
.I0(a[17]),
.I1(b[11]),
.I2(a[16]),
.I3(b[12]),
.I4(p_s0_o25_2),
.I5(1'b1));

wire p_s1_o26_4;
wire p_s1_o25_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v2 (
.O6(p_s1_o26_4),
.O5(p_s1_o25_6),
.I0(a[15]),
.I1(b[13]),
.I2(a[14]),
.I3(b[14]),
.I4(p_s0_o25_3),
.I5(1'b1));

wire p_s1_o26_5;
wire p_s1_o25_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v3 (
.O6(p_s1_o26_5),
.O5(p_s1_o25_7),
.I0(a[13]),
.I1(b[15]),
.I2(a[12]),
.I3(b[16]),
.I4(p_s0_o25_4),
.I5(1'b1));

wire p_s1_o26_6;
wire p_s1_o25_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v4 (
.O6(p_s1_o26_6),
.O5(p_s1_o25_8),
.I0(a[11]),
.I1(b[17]),
.I2(a[10]),
.I3(b[18]),
.I4(p_s0_o25_5),
.I5(1'b1));

wire p_s1_o26_7;
wire p_s1_o25_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v5 (
.O6(p_s1_o26_7),
.O5(p_s1_o25_9),
.I0(a[9]),
.I1(b[19]),
.I2(a[8]),
.I3(b[20]),
.I4(p_s0_o25_6),
.I5(1'b1));

wire p_s1_o26_8;
wire p_s1_o25_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v6 (
.O6(p_s1_o26_8),
.O5(p_s1_o25_10),
.I0(a[7]),
.I1(b[21]),
.I2(a[6]),
.I3(b[22]),
.I4(p_s0_o25_7),
.I5(1'b1));

wire p_s1_o26_9;
wire p_s1_o25_11;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v7 (
.O6(p_s1_o26_9),
.O5(p_s1_o25_11),
.I0(a[5]),
.I1(b[23]),
.I2(a[4]),
.I3(b[24]),
.I4(p_s0_o25_8),
.I5(1'b1));

wire p_s1_o26_10;
wire p_s1_o25_12;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v8 (
.O6(p_s1_o26_10),
.O5(p_s1_o25_12),
.I0(a[3]),
.I1(b[25]),
.I2(a[2]),
.I3(b[26]),
.I4(p_s0_o25_9),
.I5(1'b1));

wire p_s1_o26_11;
wire p_s1_o25_13;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o25_t81_z0_v9 (
.O6(p_s1_o26_11),
.O5(p_s1_o25_13),
.I0(a[1]),
.I1(b[27]),
.I2(a[0]),
.I3(b[28]),
.I4(p_s0_o25_10),
.I5(1'b1));

/////////STEP1----ORDER26////////////

wire p_s1_o26_12;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s1_o26_t109_z0_v0 (
.O6(p_s1_o26_12),
.O5(),
.I0(p_s0_o26_0),
.I1(p_s0_o26_1),
.I2(p_s0_o26_2),
.I3(p_s0_o26_3),
.I4(p_s0_o26_4),
.I5(p_s0_o26_5));

wire p_s1_o27_0;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s1_o26_t109_z1_v0 (
.O6(p_s1_o27_0),
.O5(),
.I0(p_s0_o26_0),
.I1(p_s0_o26_1),
.I2(p_s0_o26_2),
.I3(p_s0_o26_3),
.I4(p_s0_o26_4),
.I5(p_s0_o26_5));

wire p_s1_o28_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s1_o26_t109_z2_v0 (
.O6(p_s1_o28_0),
.O5(),
.I0(p_s0_o26_0),
.I1(p_s0_o26_1),
.I2(p_s0_o26_2),
.I3(p_s0_o26_3),
.I4(p_s0_o26_4),
.I5(p_s0_o26_5));

wire p_s1_o26_13;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s1_o26_t109_z0_v1 (
.O6(p_s1_o26_13),
.O5(),
.I0(p_s0_o26_6),
.I1(p_s0_o26_7),
.I2(p_s0_o26_8),
.I3(p_s0_o26_9),
.I4(p_s0_o26_10),
.I5(p_s0_o26_11));

wire p_s1_o27_1;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s1_o26_t109_z1_v1 (
.O6(p_s1_o27_1),
.O5(),
.I0(p_s0_o26_6),
.I1(p_s0_o26_7),
.I2(p_s0_o26_8),
.I3(p_s0_o26_9),
.I4(p_s0_o26_10),
.I5(p_s0_o26_11));

wire p_s1_o28_1;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s1_o26_t109_z2_v1 (
.O6(p_s1_o28_1),
.O5(),
.I0(p_s0_o26_6),
.I1(p_s0_o26_7),
.I2(p_s0_o26_8),
.I3(p_s0_o26_9),
.I4(p_s0_o26_10),
.I5(p_s0_o26_11));

/////////STEP1----ORDER27////////////

wire p_s1_o28_2;
wire p_s1_o27_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o27_t82_z0_v0 (
.O6(p_s1_o28_2),
.O5(p_s1_o27_2),
.I0(a[3]),
.I1(b[27]),
.I2(a[2]),
.I3(b[28]),
.I4(p_s0_o27_0),
.I5(1'b1));

wire p_s1_o28_3;
wire p_s1_o27_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o27_t82_z0_v1 (
.O6(p_s1_o28_3),
.O5(p_s1_o27_3),
.I0(a[1]),
.I1(b[29]),
.I2(a[0]),
.I3(b[30]),
.I4(p_s0_o27_1),
.I5(1'b1));

wire p_s1_o27_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o27_t113_z0_v0 (
.O6(p_s1_o27_4),
.O5(),
.I0(p_s0_o27_2),
.I1(p_s0_o27_3),
.I2(p_s0_o27_4),
.I3(p_s0_o27_5),
.I4(p_s0_o27_6),
.I5(p_s0_o28_0));

wire p_s1_o28_4;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o27_t113_z1_v0 (
.O6(p_s1_o28_4),
.O5(),
.I0(p_s0_o27_2),
.I1(p_s0_o27_3),
.I2(p_s0_o27_4),
.I3(p_s0_o27_5),
.I4(p_s0_o27_6),
.I5(p_s0_o28_0));

wire p_s1_o29_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o27_t113_z2_v0 (
.O6(p_s1_o29_0),
.O5(),
.I0(p_s0_o27_2),
.I1(p_s0_o27_3),
.I2(p_s0_o27_4),
.I3(p_s0_o27_5),
.I4(p_s0_o27_6),
.I5(p_s0_o28_0));

wire p_s1_o27_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o27_t113_z0_v1 (
.O6(p_s1_o27_5),
.O5(),
.I0(p_s0_o27_7),
.I1(p_s0_o27_8),
.I2(p_s0_o27_9),
.I3(p_s0_o27_10),
.I4(p_s0_o27_11),
.I5(p_s0_o28_1));

wire p_s1_o28_5;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o27_t113_z1_v1 (
.O6(p_s1_o28_5),
.O5(),
.I0(p_s0_o27_7),
.I1(p_s0_o27_8),
.I2(p_s0_o27_9),
.I3(p_s0_o27_10),
.I4(p_s0_o27_11),
.I5(p_s0_o28_1));

wire p_s1_o29_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o27_t113_z2_v1 (
.O6(p_s1_o29_1),
.O5(),
.I0(p_s0_o27_7),
.I1(p_s0_o27_8),
.I2(p_s0_o27_9),
.I3(p_s0_o27_10),
.I4(p_s0_o27_11),
.I5(p_s0_o28_1));

wire p_s1_o27_6;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o27_t113_z0_v2 (
.O6(p_s1_o27_6),
.O5(),
.I0(p_s0_o27_12),
.I1(p_s0_o27_13),
.I2(p_s0_o27_14),
.I3(p_s0_o27_15),
.I4(p_s0_o27_16),
.I5(p_s0_o28_2));

wire p_s1_o28_6;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o27_t113_z1_v2 (
.O6(p_s1_o28_6),
.O5(),
.I0(p_s0_o27_12),
.I1(p_s0_o27_13),
.I2(p_s0_o27_14),
.I3(p_s0_o27_15),
.I4(p_s0_o27_16),
.I5(p_s0_o28_2));

wire p_s1_o29_2;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o27_t113_z2_v2 (
.O6(p_s1_o29_2),
.O5(),
.I0(p_s0_o27_12),
.I1(p_s0_o27_13),
.I2(p_s0_o27_14),
.I3(p_s0_o27_15),
.I4(p_s0_o27_16),
.I5(p_s0_o28_2));

/////////STEP1----ORDER28////////////

wire p_s1_o29_3;
wire p_s1_o28_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o28_t83_z0_v0 (
.O6(p_s1_o29_3),
.O5(p_s1_o28_7),
.I0(a[1]),
.I1(b[30]),
.I2(a[0]),
.I3(b[31]),
.I4(p_s0_o28_3),
.I5(1'b1));

wire p_s1_o28_8;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o28_t114_z0_v0 (
.O6(p_s1_o28_8),
.O5(),
.I0(p_s0_o28_4),
.I1(p_s0_o28_5),
.I2(p_s0_o28_6),
.I3(p_s0_o28_7),
.I4(p_s0_o28_8),
.I5(p_s0_o29_0));

wire p_s1_o29_4;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o28_t114_z1_v0 (
.O6(p_s1_o29_4),
.O5(),
.I0(p_s0_o28_4),
.I1(p_s0_o28_5),
.I2(p_s0_o28_6),
.I3(p_s0_o28_7),
.I4(p_s0_o28_8),
.I5(p_s0_o29_0));

wire p_s1_o30_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o28_t114_z2_v0 (
.O6(p_s1_o30_0),
.O5(),
.I0(p_s0_o28_4),
.I1(p_s0_o28_5),
.I2(p_s0_o28_6),
.I3(p_s0_o28_7),
.I4(p_s0_o28_8),
.I5(p_s0_o29_0));

wire p_s1_o28_9;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o28_t114_z0_v1 (
.O6(p_s1_o28_9),
.O5(),
.I0(p_s0_o28_9),
.I1(p_s0_o28_10),
.I2(p_s0_o28_11),
.I3(p_s0_o28_12),
.I4(p_s0_o28_13),
.I5(p_s0_o29_1));

wire p_s1_o29_5;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o28_t114_z1_v1 (
.O6(p_s1_o29_5),
.O5(),
.I0(p_s0_o28_9),
.I1(p_s0_o28_10),
.I2(p_s0_o28_11),
.I3(p_s0_o28_12),
.I4(p_s0_o28_13),
.I5(p_s0_o29_1));

wire p_s1_o30_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o28_t114_z2_v1 (
.O6(p_s1_o30_1),
.O5(),
.I0(p_s0_o28_9),
.I1(p_s0_o28_10),
.I2(p_s0_o28_11),
.I3(p_s0_o28_12),
.I4(p_s0_o28_13),
.I5(p_s0_o29_1));

wire p_s1_o28_10;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o28_t114_z0_v2 (
.O6(p_s1_o28_10),
.O5(),
.I0(p_s0_o28_14),
.I1(p_s0_o28_15),
.I2(p_s0_o28_16),
.I3(p_s0_o28_17),
.I4(p_s0_o28_18),
.I5(p_s0_o29_2));

wire p_s1_o29_6;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o28_t114_z1_v2 (
.O6(p_s1_o29_6),
.O5(),
.I0(p_s0_o28_14),
.I1(p_s0_o28_15),
.I2(p_s0_o28_16),
.I3(p_s0_o28_17),
.I4(p_s0_o28_18),
.I5(p_s0_o29_2));

wire p_s1_o30_2;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o28_t114_z2_v2 (
.O6(p_s1_o30_2),
.O5(),
.I0(p_s0_o28_14),
.I1(p_s0_o28_15),
.I2(p_s0_o28_16),
.I3(p_s0_o28_17),
.I4(p_s0_o28_18),
.I5(p_s0_o29_2));

/////////STEP1----ORDER29////////////

wire p_s1_o30_3;
wire p_s1_o29_7;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o29_t52_z0_v0 (
.O6(p_s1_o30_3),
.O5(p_s1_o29_7),
.I0(a[1]),
.I1(b[31]),
.I2(p_s0_o29_3),
.I3(p_s0_o29_4),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o29_8;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o29_t115_z0_v0 (
.O6(p_s1_o29_8),
.O5(),
.I0(p_s0_o29_5),
.I1(p_s0_o29_6),
.I2(p_s0_o29_7),
.I3(p_s0_o29_8),
.I4(p_s0_o29_9),
.I5(p_s0_o30_0));

wire p_s1_o30_4;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o29_t115_z1_v0 (
.O6(p_s1_o30_4),
.O5(),
.I0(p_s0_o29_5),
.I1(p_s0_o29_6),
.I2(p_s0_o29_7),
.I3(p_s0_o29_8),
.I4(p_s0_o29_9),
.I5(p_s0_o30_0));

wire p_s1_o31_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o29_t115_z2_v0 (
.O6(p_s1_o31_0),
.O5(),
.I0(p_s0_o29_5),
.I1(p_s0_o29_6),
.I2(p_s0_o29_7),
.I3(p_s0_o29_8),
.I4(p_s0_o29_9),
.I5(p_s0_o30_0));

wire p_s1_o29_9;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o29_t115_z0_v1 (
.O6(p_s1_o29_9),
.O5(),
.I0(p_s0_o29_10),
.I1(p_s0_o29_11),
.I2(p_s0_o29_12),
.I3(p_s0_o29_13),
.I4(p_s0_o29_14),
.I5(p_s0_o30_1));

wire p_s1_o30_5;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o29_t115_z1_v1 (
.O6(p_s1_o30_5),
.O5(),
.I0(p_s0_o29_10),
.I1(p_s0_o29_11),
.I2(p_s0_o29_12),
.I3(p_s0_o29_13),
.I4(p_s0_o29_14),
.I5(p_s0_o30_1));

wire p_s1_o31_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o29_t115_z2_v1 (
.O6(p_s1_o31_1),
.O5(),
.I0(p_s0_o29_10),
.I1(p_s0_o29_11),
.I2(p_s0_o29_12),
.I3(p_s0_o29_13),
.I4(p_s0_o29_14),
.I5(p_s0_o30_1));

wire p_s1_o29_10;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o29_t115_z0_v2 (
.O6(p_s1_o29_10),
.O5(),
.I0(p_s0_o29_15),
.I1(p_s0_o29_16),
.I2(p_s0_o29_17),
.I3(p_s0_o29_18),
.I4(p_s0_o29_19),
.I5(p_s0_o30_2));

wire p_s1_o30_6;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o29_t115_z1_v2 (
.O6(p_s1_o30_6),
.O5(),
.I0(p_s0_o29_15),
.I1(p_s0_o29_16),
.I2(p_s0_o29_17),
.I3(p_s0_o29_18),
.I4(p_s0_o29_19),
.I5(p_s0_o30_2));

wire p_s1_o31_2;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o29_t115_z2_v2 (
.O6(p_s1_o31_2),
.O5(),
.I0(p_s0_o29_15),
.I1(p_s0_o29_16),
.I2(p_s0_o29_17),
.I3(p_s0_o29_18),
.I4(p_s0_o29_19),
.I5(p_s0_o30_2));

/////////STEP1----ORDER30////////////

wire p_s1_o31_3;
wire p_s1_o30_7;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s1_o30_t48_z0_v0 (
.O6(p_s1_o31_3),
.O5(p_s1_o30_7),
.I0(p_s0_o30_3),
.I1(p_s0_o30_4),
.I2(p_s0_o30_5),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o31_4;
wire p_s1_o30_8;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o30_t53_z0_v0 (
.O6(p_s1_o31_4),
.O5(p_s1_o30_8),
.I0(a[4]),
.I1(b[29]),
.I2(p_s0_o30_6),
.I3(p_s0_o30_7),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o31_5;
wire p_s1_o30_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o30_t84_z0_v0 (
.O6(p_s1_o31_5),
.O5(p_s1_o30_9),
.I0(a[3]),
.I1(b[30]),
.I2(a[2]),
.I3(b[31]),
.I4(p_s0_o30_8),
.I5(1'b1));

wire p_s1_o30_10;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o30_t116_z0_v0 (
.O6(p_s1_o30_10),
.O5(),
.I0(p_s0_o30_9),
.I1(p_s0_o30_10),
.I2(p_s0_o30_11),
.I3(p_s0_o30_12),
.I4(p_s0_o30_13),
.I5(p_s0_o31_0));

wire p_s1_o31_6;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o30_t116_z1_v0 (
.O6(p_s1_o31_6),
.O5(),
.I0(p_s0_o30_9),
.I1(p_s0_o30_10),
.I2(p_s0_o30_11),
.I3(p_s0_o30_12),
.I4(p_s0_o30_13),
.I5(p_s0_o31_0));

wire p_s1_o32_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o30_t116_z2_v0 (
.O6(p_s1_o32_0),
.O5(),
.I0(p_s0_o30_9),
.I1(p_s0_o30_10),
.I2(p_s0_o30_11),
.I3(p_s0_o30_12),
.I4(p_s0_o30_13),
.I5(p_s0_o31_0));

wire p_s1_o30_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o30_t116_z0_v1 (
.O6(p_s1_o30_11),
.O5(),
.I0(p_s0_o30_14),
.I1(p_s0_o30_15),
.I2(p_s0_o30_16),
.I3(p_s0_o30_17),
.I4(p_s0_o30_18),
.I5(p_s0_o31_1));

wire p_s1_o31_7;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o30_t116_z1_v1 (
.O6(p_s1_o31_7),
.O5(),
.I0(p_s0_o30_14),
.I1(p_s0_o30_15),
.I2(p_s0_o30_16),
.I3(p_s0_o30_17),
.I4(p_s0_o30_18),
.I5(p_s0_o31_1));

wire p_s1_o32_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o30_t116_z2_v1 (
.O6(p_s1_o32_1),
.O5(),
.I0(p_s0_o30_14),
.I1(p_s0_o30_15),
.I2(p_s0_o30_16),
.I3(p_s0_o30_17),
.I4(p_s0_o30_18),
.I5(p_s0_o31_1));

/////////STEP1----ORDER31////////////

wire p_s1_o32_2;
wire p_s1_o31_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o31_t85_z0_v0 (
.O6(p_s1_o32_2),
.O5(p_s1_o31_8),
.I0(a[4]),
.I1(b[30]),
.I2(a[3]),
.I3(b[31]),
.I4(p_s0_o31_2),
.I5(1'b1));

wire p_s1_o31_9;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o31_t117_z0_v0 (
.O6(p_s1_o31_9),
.O5(),
.I0(p_s0_o31_3),
.I1(p_s0_o31_4),
.I2(p_s0_o31_5),
.I3(p_s0_o31_6),
.I4(p_s0_o31_7),
.I5(p_s0_o32_0));

wire p_s1_o32_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o31_t117_z1_v0 (
.O6(p_s1_o32_3),
.O5(),
.I0(p_s0_o31_3),
.I1(p_s0_o31_4),
.I2(p_s0_o31_5),
.I3(p_s0_o31_6),
.I4(p_s0_o31_7),
.I5(p_s0_o32_0));

wire p_s1_o33_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o31_t117_z2_v0 (
.O6(p_s1_o33_0),
.O5(),
.I0(p_s0_o31_3),
.I1(p_s0_o31_4),
.I2(p_s0_o31_5),
.I3(p_s0_o31_6),
.I4(p_s0_o31_7),
.I5(p_s0_o32_0));

wire p_s1_o31_10;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o31_t117_z0_v1 (
.O6(p_s1_o31_10),
.O5(),
.I0(p_s0_o31_8),
.I1(p_s0_o31_9),
.I2(p_s0_o31_10),
.I3(p_s0_o31_11),
.I4(p_s0_o31_12),
.I5(p_s0_o32_1));

wire p_s1_o32_4;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o31_t117_z1_v1 (
.O6(p_s1_o32_4),
.O5(),
.I0(p_s0_o31_8),
.I1(p_s0_o31_9),
.I2(p_s0_o31_10),
.I3(p_s0_o31_11),
.I4(p_s0_o31_12),
.I5(p_s0_o32_1));

wire p_s1_o33_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o31_t117_z2_v1 (
.O6(p_s1_o33_1),
.O5(),
.I0(p_s0_o31_8),
.I1(p_s0_o31_9),
.I2(p_s0_o31_10),
.I3(p_s0_o31_11),
.I4(p_s0_o31_12),
.I5(p_s0_o32_1));

wire p_s1_o31_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o31_t117_z0_v2 (
.O6(p_s1_o31_11),
.O5(),
.I0(p_s0_o31_13),
.I1(p_s0_o31_14),
.I2(p_s0_o31_15),
.I3(p_s0_o31_16),
.I4(p_s0_o31_17),
.I5(p_s0_o32_2));

wire p_s1_o32_5;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o31_t117_z1_v2 (
.O6(p_s1_o32_5),
.O5(),
.I0(p_s0_o31_13),
.I1(p_s0_o31_14),
.I2(p_s0_o31_15),
.I3(p_s0_o31_16),
.I4(p_s0_o31_17),
.I5(p_s0_o32_2));

wire p_s1_o33_2;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o31_t117_z2_v2 (
.O6(p_s1_o33_2),
.O5(),
.I0(p_s0_o31_13),
.I1(p_s0_o31_14),
.I2(p_s0_o31_15),
.I3(p_s0_o31_16),
.I4(p_s0_o31_17),
.I5(p_s0_o32_2));

/////////STEP1----ORDER32////////////

wire p_s1_o33_3;
wire p_s1_o32_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o32_t86_z0_v0 (
.O6(p_s1_o33_3),
.O5(p_s1_o32_6),
.I0(a[7]),
.I1(b[28]),
.I2(a[6]),
.I3(b[29]),
.I4(p_s0_o32_3),
.I5(1'b1));

wire p_s1_o33_4;
wire p_s1_o32_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o32_t86_z0_v1 (
.O6(p_s1_o33_4),
.O5(p_s1_o32_7),
.I0(a[5]),
.I1(b[30]),
.I2(a[4]),
.I3(b[31]),
.I4(p_s0_o32_4),
.I5(1'b1));

wire p_s1_o32_8;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o32_t118_z0_v0 (
.O6(p_s1_o32_8),
.O5(),
.I0(p_s0_o32_5),
.I1(p_s0_o32_6),
.I2(p_s0_o32_7),
.I3(p_s0_o32_8),
.I4(p_s0_o32_9),
.I5(p_s0_o33_0));

wire p_s1_o33_5;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o32_t118_z1_v0 (
.O6(p_s1_o33_5),
.O5(),
.I0(p_s0_o32_5),
.I1(p_s0_o32_6),
.I2(p_s0_o32_7),
.I3(p_s0_o32_8),
.I4(p_s0_o32_9),
.I5(p_s0_o33_0));

wire p_s1_o34_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o32_t118_z2_v0 (
.O6(p_s1_o34_0),
.O5(),
.I0(p_s0_o32_5),
.I1(p_s0_o32_6),
.I2(p_s0_o32_7),
.I3(p_s0_o32_8),
.I4(p_s0_o32_9),
.I5(p_s0_o33_0));

wire p_s1_o32_9;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o32_t118_z0_v1 (
.O6(p_s1_o32_9),
.O5(),
.I0(p_s0_o32_10),
.I1(p_s0_o32_11),
.I2(p_s0_o32_12),
.I3(p_s0_o32_13),
.I4(p_s0_o32_14),
.I5(p_s0_o33_1));

wire p_s1_o33_6;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o32_t118_z1_v1 (
.O6(p_s1_o33_6),
.O5(),
.I0(p_s0_o32_10),
.I1(p_s0_o32_11),
.I2(p_s0_o32_12),
.I3(p_s0_o32_13),
.I4(p_s0_o32_14),
.I5(p_s0_o33_1));

wire p_s1_o34_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o32_t118_z2_v1 (
.O6(p_s1_o34_1),
.O5(),
.I0(p_s0_o32_10),
.I1(p_s0_o32_11),
.I2(p_s0_o32_12),
.I3(p_s0_o32_13),
.I4(p_s0_o32_14),
.I5(p_s0_o33_1));

/////////STEP1----ORDER33////////////

wire p_s1_o34_2;
wire p_s1_o33_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o33_t87_z0_v0 (
.O6(p_s1_o34_2),
.O5(p_s1_o33_7),
.I0(a[10]),
.I1(b[26]),
.I2(a[9]),
.I3(b[27]),
.I4(p_s0_o33_2),
.I5(1'b1));

wire p_s1_o34_3;
wire p_s1_o33_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o33_t87_z0_v1 (
.O6(p_s1_o34_3),
.O5(p_s1_o33_8),
.I0(a[8]),
.I1(b[28]),
.I2(a[7]),
.I3(b[29]),
.I4(p_s0_o33_3),
.I5(1'b1));

wire p_s1_o34_4;
wire p_s1_o33_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o33_t87_z0_v2 (
.O6(p_s1_o34_4),
.O5(p_s1_o33_9),
.I0(a[6]),
.I1(b[30]),
.I2(a[5]),
.I3(b[31]),
.I4(p_s0_o33_4),
.I5(1'b1));

wire p_s1_o33_10;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o33_t119_z0_v0 (
.O6(p_s1_o33_10),
.O5(),
.I0(p_s0_o33_5),
.I1(p_s0_o33_6),
.I2(p_s0_o33_7),
.I3(p_s0_o33_8),
.I4(p_s0_o33_9),
.I5(p_s0_o34_0));

wire p_s1_o34_5;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o33_t119_z1_v0 (
.O6(p_s1_o34_5),
.O5(),
.I0(p_s0_o33_5),
.I1(p_s0_o33_6),
.I2(p_s0_o33_7),
.I3(p_s0_o33_8),
.I4(p_s0_o33_9),
.I5(p_s0_o34_0));

wire p_s1_o35_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o33_t119_z2_v0 (
.O6(p_s1_o35_0),
.O5(),
.I0(p_s0_o33_5),
.I1(p_s0_o33_6),
.I2(p_s0_o33_7),
.I3(p_s0_o33_8),
.I4(p_s0_o33_9),
.I5(p_s0_o34_0));

wire p_s1_o33_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o33_t119_z0_v1 (
.O6(p_s1_o33_11),
.O5(),
.I0(p_s0_o33_10),
.I1(p_s0_o33_11),
.I2(p_s0_o33_12),
.I3(p_s0_o33_13),
.I4(p_s0_o33_14),
.I5(p_s0_o34_1));

wire p_s1_o34_6;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o33_t119_z1_v1 (
.O6(p_s1_o34_6),
.O5(),
.I0(p_s0_o33_10),
.I1(p_s0_o33_11),
.I2(p_s0_o33_12),
.I3(p_s0_o33_13),
.I4(p_s0_o33_14),
.I5(p_s0_o34_1));

wire p_s1_o35_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o33_t119_z2_v1 (
.O6(p_s1_o35_1),
.O5(),
.I0(p_s0_o33_10),
.I1(p_s0_o33_11),
.I2(p_s0_o33_12),
.I3(p_s0_o33_13),
.I4(p_s0_o33_14),
.I5(p_s0_o34_1));

/////////STEP1----ORDER34////////////

wire p_s1_o35_2;
wire p_s1_o34_7;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s1_o34_t49_z0_v0 (
.O6(p_s1_o35_2),
.O5(p_s1_o34_7),
.I0(p_s0_o34_2),
.I1(p_s0_o34_3),
.I2(p_s0_o34_4),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o35_3;
wire p_s1_o34_8;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o34_t54_z0_v0 (
.O6(p_s1_o35_3),
.O5(p_s1_o34_8),
.I0(a[10]),
.I1(b[27]),
.I2(p_s0_o34_5),
.I3(p_s0_o34_6),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o35_4;
wire p_s1_o34_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o34_t88_z0_v0 (
.O6(p_s1_o35_4),
.O5(p_s1_o34_9),
.I0(a[9]),
.I1(b[28]),
.I2(a[8]),
.I3(b[29]),
.I4(p_s0_o34_7),
.I5(1'b1));

wire p_s1_o35_5;
wire p_s1_o34_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o34_t88_z0_v1 (
.O6(p_s1_o35_5),
.O5(p_s1_o34_10),
.I0(a[7]),
.I1(b[30]),
.I2(a[6]),
.I3(b[31]),
.I4(p_s0_o34_8),
.I5(1'b1));

wire p_s1_o34_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o34_t120_z0_v0 (
.O6(p_s1_o34_11),
.O5(),
.I0(p_s0_o34_9),
.I1(p_s0_o34_10),
.I2(p_s0_o34_11),
.I3(p_s0_o34_12),
.I4(p_s0_o34_13),
.I5(p_s0_o35_0));

wire p_s1_o35_6;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o34_t120_z1_v0 (
.O6(p_s1_o35_6),
.O5(),
.I0(p_s0_o34_9),
.I1(p_s0_o34_10),
.I2(p_s0_o34_11),
.I3(p_s0_o34_12),
.I4(p_s0_o34_13),
.I5(p_s0_o35_0));

wire p_s1_o36_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o34_t120_z2_v0 (
.O6(p_s1_o36_0),
.O5(),
.I0(p_s0_o34_9),
.I1(p_s0_o34_10),
.I2(p_s0_o34_11),
.I3(p_s0_o34_12),
.I4(p_s0_o34_13),
.I5(p_s0_o35_0));

/////////STEP1----ORDER35////////////

wire p_s1_o36_1;
wire p_s1_o35_7;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s1_o35_t50_z0_v0 (
.O6(p_s1_o36_1),
.O5(p_s1_o35_7),
.I0(p_s0_o35_1),
.I1(p_s0_o35_2),
.I2(p_s0_o35_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o36_2;
wire p_s1_o35_8;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s1_o35_t50_z0_v1 (
.O6(p_s1_o36_2),
.O5(p_s1_o35_8),
.I0(p_s0_o35_4),
.I1(p_s0_o35_5),
.I2(p_s0_o35_6),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o36_3;
wire p_s1_o35_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o35_t89_z0_v0 (
.O6(p_s1_o36_3),
.O5(p_s1_o35_9),
.I0(a[10]),
.I1(b[28]),
.I2(a[9]),
.I3(b[29]),
.I4(p_s0_o35_7),
.I5(1'b1));

wire p_s1_o36_4;
wire p_s1_o35_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o35_t89_z0_v1 (
.O6(p_s1_o36_4),
.O5(p_s1_o35_10),
.I0(a[8]),
.I1(b[30]),
.I2(a[7]),
.I3(b[31]),
.I4(p_s0_o35_8),
.I5(1'b1));

wire p_s1_o35_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o35_t121_z0_v0 (
.O6(p_s1_o35_11),
.O5(),
.I0(p_s0_o35_9),
.I1(p_s0_o35_10),
.I2(p_s0_o35_11),
.I3(p_s0_o35_12),
.I4(p_s0_o35_13),
.I5(p_s0_o36_0));

wire p_s1_o36_5;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o35_t121_z1_v0 (
.O6(p_s1_o36_5),
.O5(),
.I0(p_s0_o35_9),
.I1(p_s0_o35_10),
.I2(p_s0_o35_11),
.I3(p_s0_o35_12),
.I4(p_s0_o35_13),
.I5(p_s0_o36_0));

wire p_s1_o37_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o35_t121_z2_v0 (
.O6(p_s1_o37_0),
.O5(),
.I0(p_s0_o35_9),
.I1(p_s0_o35_10),
.I2(p_s0_o35_11),
.I3(p_s0_o35_12),
.I4(p_s0_o35_13),
.I5(p_s0_o36_0));

/////////STEP1----ORDER36////////////

wire p_s1_o37_1;
wire p_s1_o36_6;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o36_t55_z0_v0 (
.O6(p_s1_o37_1),
.O5(p_s1_o36_6),
.I0(a[16]),
.I1(b[23]),
.I2(p_s0_o36_1),
.I3(p_s0_o36_2),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o37_2;
wire p_s1_o36_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o36_t90_z0_v0 (
.O6(p_s1_o37_2),
.O5(p_s1_o36_7),
.I0(a[15]),
.I1(b[24]),
.I2(a[14]),
.I3(b[25]),
.I4(p_s0_o36_3),
.I5(1'b1));

wire p_s1_o37_3;
wire p_s1_o36_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o36_t90_z0_v1 (
.O6(p_s1_o37_3),
.O5(p_s1_o36_8),
.I0(a[13]),
.I1(b[26]),
.I2(a[12]),
.I3(b[27]),
.I4(p_s0_o36_4),
.I5(1'b1));

wire p_s1_o37_4;
wire p_s1_o36_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o36_t90_z0_v2 (
.O6(p_s1_o37_4),
.O5(p_s1_o36_9),
.I0(a[11]),
.I1(b[28]),
.I2(a[10]),
.I3(b[29]),
.I4(p_s0_o36_5),
.I5(1'b1));

wire p_s1_o37_5;
wire p_s1_o36_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o36_t90_z0_v3 (
.O6(p_s1_o37_5),
.O5(p_s1_o36_10),
.I0(a[9]),
.I1(b[30]),
.I2(a[8]),
.I3(b[31]),
.I4(p_s0_o36_6),
.I5(1'b1));

wire p_s1_o36_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o36_t122_z0_v0 (
.O6(p_s1_o36_11),
.O5(),
.I0(p_s0_o36_7),
.I1(p_s0_o36_8),
.I2(p_s0_o36_9),
.I3(p_s0_o36_10),
.I4(p_s0_o36_11),
.I5(p_s0_o37_0));

wire p_s1_o37_6;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o36_t122_z1_v0 (
.O6(p_s1_o37_6),
.O5(),
.I0(p_s0_o36_7),
.I1(p_s0_o36_8),
.I2(p_s0_o36_9),
.I3(p_s0_o36_10),
.I4(p_s0_o36_11),
.I5(p_s0_o37_0));

wire p_s1_o38_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o36_t122_z2_v0 (
.O6(p_s1_o38_0),
.O5(),
.I0(p_s0_o36_7),
.I1(p_s0_o36_8),
.I2(p_s0_o36_9),
.I3(p_s0_o36_10),
.I4(p_s0_o36_11),
.I5(p_s0_o37_0));

/////////STEP1----ORDER37////////////

wire p_s1_o38_1;
wire p_s1_o37_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o37_t91_z0_v0 (
.O6(p_s1_o38_1),
.O5(p_s1_o37_7),
.I0(a[16]),
.I1(b[24]),
.I2(a[15]),
.I3(b[25]),
.I4(p_s0_o37_1),
.I5(1'b1));

wire p_s1_o38_2;
wire p_s1_o37_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o37_t91_z0_v1 (
.O6(p_s1_o38_2),
.O5(p_s1_o37_8),
.I0(a[14]),
.I1(b[26]),
.I2(a[13]),
.I3(b[27]),
.I4(p_s0_o37_2),
.I5(1'b1));

wire p_s1_o38_3;
wire p_s1_o37_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o37_t91_z0_v2 (
.O6(p_s1_o38_3),
.O5(p_s1_o37_9),
.I0(a[12]),
.I1(b[28]),
.I2(a[11]),
.I3(b[29]),
.I4(p_s0_o37_3),
.I5(1'b1));

wire p_s1_o38_4;
wire p_s1_o37_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o37_t91_z0_v3 (
.O6(p_s1_o38_4),
.O5(p_s1_o37_10),
.I0(a[10]),
.I1(b[30]),
.I2(a[9]),
.I3(b[31]),
.I4(p_s0_o37_4),
.I5(1'b1));

wire p_s1_o37_11;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s1_o37_t123_z0_v0 (
.O6(p_s1_o37_11),
.O5(),
.I0(p_s0_o37_5),
.I1(p_s0_o37_6),
.I2(p_s0_o37_7),
.I3(p_s0_o37_8),
.I4(p_s0_o37_9),
.I5(p_s0_o38_0));

wire p_s1_o38_5;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s1_o37_t123_z1_v0 (
.O6(p_s1_o38_5),
.O5(),
.I0(p_s0_o37_5),
.I1(p_s0_o37_6),
.I2(p_s0_o37_7),
.I3(p_s0_o37_8),
.I4(p_s0_o37_9),
.I5(p_s0_o38_0));

wire p_s1_o39_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s1_o37_t123_z2_v0 (
.O6(p_s1_o39_0),
.O5(),
.I0(p_s0_o37_5),
.I1(p_s0_o37_6),
.I2(p_s0_o37_7),
.I3(p_s0_o37_8),
.I4(p_s0_o37_9),
.I5(p_s0_o38_0));

/////////STEP1----ORDER38////////////

wire p_s1_o39_1;
wire p_s1_o38_6;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o38_t56_z0_v0 (
.O6(p_s1_o39_1),
.O5(p_s1_o38_6),
.I0(a[19]),
.I1(b[22]),
.I2(p_s0_o38_1),
.I3(p_s0_o38_2),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o39_2;
wire p_s1_o38_7;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o38_t56_z0_v1 (
.O6(p_s1_o39_2),
.O5(p_s1_o38_7),
.I0(a[18]),
.I1(b[23]),
.I2(p_s0_o38_3),
.I3(p_s0_o38_4),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o39_3;
wire p_s1_o38_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o38_t92_z0_v0 (
.O6(p_s1_o39_3),
.O5(p_s1_o38_8),
.I0(a[17]),
.I1(b[24]),
.I2(a[16]),
.I3(b[25]),
.I4(p_s0_o38_5),
.I5(1'b1));

wire p_s1_o39_4;
wire p_s1_o38_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o38_t92_z0_v1 (
.O6(p_s1_o39_4),
.O5(p_s1_o38_9),
.I0(a[15]),
.I1(b[26]),
.I2(a[14]),
.I3(b[27]),
.I4(p_s0_o38_6),
.I5(1'b1));

wire p_s1_o39_5;
wire p_s1_o38_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o38_t92_z0_v2 (
.O6(p_s1_o39_5),
.O5(p_s1_o38_10),
.I0(a[13]),
.I1(b[28]),
.I2(a[12]),
.I3(b[29]),
.I4(p_s0_o38_7),
.I5(1'b1));

wire p_s1_o39_6;
wire p_s1_o38_11;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o38_t92_z0_v3 (
.O6(p_s1_o39_6),
.O5(p_s1_o38_11),
.I0(a[11]),
.I1(b[30]),
.I2(a[10]),
.I3(b[31]),
.I4(p_s0_o38_8),
.I5(1'b1));

/////////STEP1----ORDER39////////////

wire p_s1_o40_0;
wire p_s1_o39_7;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o39_t57_z0_v0 (
.O6(p_s1_o40_0),
.O5(p_s1_o39_7),
.I0(a[16]),
.I1(b[26]),
.I2(p_s0_o39_0),
.I3(p_s0_o39_1),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o40_1;
wire p_s1_o39_8;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o39_t57_z0_v1 (
.O6(p_s1_o40_1),
.O5(p_s1_o39_8),
.I0(a[15]),
.I1(b[27]),
.I2(p_s0_o39_2),
.I3(p_s0_o39_3),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o40_2;
wire p_s1_o39_9;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o39_t57_z0_v2 (
.O6(p_s1_o40_2),
.O5(p_s1_o39_9),
.I0(a[14]),
.I1(b[28]),
.I2(p_s0_o39_4),
.I3(p_s0_o39_5),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o40_3;
wire p_s1_o39_10;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o39_t57_z0_v3 (
.O6(p_s1_o40_3),
.O5(p_s1_o39_10),
.I0(a[13]),
.I1(b[29]),
.I2(p_s0_o39_6),
.I3(p_s0_o39_7),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o40_4;
wire p_s1_o39_11;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o39_t93_z0_v0 (
.O6(p_s1_o40_4),
.O5(p_s1_o39_11),
.I0(a[12]),
.I1(b[30]),
.I2(a[11]),
.I3(b[31]),
.I4(p_s0_o39_8),
.I5(1'b1));

/////////STEP1----ORDER40////////////

wire p_s1_o41_0;
wire p_s1_o40_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o40_t94_z0_v0 (
.O6(p_s1_o41_0),
.O5(p_s1_o40_5),
.I0(a[25]),
.I1(b[18]),
.I2(a[24]),
.I3(b[19]),
.I4(p_s0_o40_0),
.I5(1'b1));

wire p_s1_o41_1;
wire p_s1_o40_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o40_t94_z0_v1 (
.O6(p_s1_o41_1),
.O5(p_s1_o40_6),
.I0(a[23]),
.I1(b[20]),
.I2(a[22]),
.I3(b[21]),
.I4(p_s0_o40_1),
.I5(1'b1));

wire p_s1_o41_2;
wire p_s1_o40_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o40_t94_z0_v2 (
.O6(p_s1_o41_2),
.O5(p_s1_o40_7),
.I0(a[21]),
.I1(b[22]),
.I2(a[20]),
.I3(b[23]),
.I4(p_s0_o40_2),
.I5(1'b1));

wire p_s1_o41_3;
wire p_s1_o40_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o40_t94_z0_v3 (
.O6(p_s1_o41_3),
.O5(p_s1_o40_8),
.I0(a[19]),
.I1(b[24]),
.I2(a[18]),
.I3(b[25]),
.I4(p_s0_o40_3),
.I5(1'b1));

wire p_s1_o41_4;
wire p_s1_o40_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o40_t94_z0_v4 (
.O6(p_s1_o41_4),
.O5(p_s1_o40_9),
.I0(a[17]),
.I1(b[26]),
.I2(a[16]),
.I3(b[27]),
.I4(p_s0_o40_4),
.I5(1'b1));

wire p_s1_o41_5;
wire p_s1_o40_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o40_t94_z0_v5 (
.O6(p_s1_o41_5),
.O5(p_s1_o40_10),
.I0(a[15]),
.I1(b[28]),
.I2(a[14]),
.I3(b[29]),
.I4(p_s0_o40_5),
.I5(1'b1));

wire p_s1_o41_6;
wire p_s1_o40_11;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o40_t94_z0_v6 (
.O6(p_s1_o41_6),
.O5(p_s1_o40_11),
.I0(a[13]),
.I1(b[30]),
.I2(a[12]),
.I3(b[31]),
.I4(p_s0_o40_6),
.I5(1'b1));

/////////STEP1----ORDER41////////////

wire p_s1_o42_0;
wire p_s1_o41_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o41_t95_z0_v0 (
.O6(p_s1_o42_0),
.O5(p_s1_o41_7),
.I0(a[22]),
.I1(b[22]),
.I2(a[21]),
.I3(b[23]),
.I4(p_s0_o41_0),
.I5(1'b1));

wire p_s1_o42_1;
wire p_s1_o41_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o41_t95_z0_v1 (
.O6(p_s1_o42_1),
.O5(p_s1_o41_8),
.I0(a[20]),
.I1(b[24]),
.I2(a[19]),
.I3(b[25]),
.I4(p_s0_o41_1),
.I5(1'b1));

wire p_s1_o42_2;
wire p_s1_o41_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o41_t95_z0_v2 (
.O6(p_s1_o42_2),
.O5(p_s1_o41_9),
.I0(a[18]),
.I1(b[26]),
.I2(a[17]),
.I3(b[27]),
.I4(p_s0_o41_2),
.I5(1'b1));

wire p_s1_o42_3;
wire p_s1_o41_10;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o41_t95_z0_v3 (
.O6(p_s1_o42_3),
.O5(p_s1_o41_10),
.I0(a[16]),
.I1(b[28]),
.I2(a[15]),
.I3(b[29]),
.I4(p_s0_o41_3),
.I5(1'b1));

wire p_s1_o42_4;
wire p_s1_o41_11;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o41_t95_z0_v4 (
.O6(p_s1_o42_4),
.O5(p_s1_o41_11),
.I0(a[14]),
.I1(b[30]),
.I2(a[13]),
.I3(b[31]),
.I4(p_s0_o41_4),
.I5(1'b1));

/////////STEP1----ORDER42////////////

wire p_s1_o43_0;
wire p_s1_o42_5;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o42_t58_z0_v0 (
.O6(p_s1_o43_0),
.O5(p_s1_o42_5),
.I0(a[22]),
.I1(b[23]),
.I2(p_s0_o42_0),
.I3(p_s0_o42_1),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o43_1;
wire p_s1_o42_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o42_t96_z0_v0 (
.O6(p_s1_o43_1),
.O5(p_s1_o42_6),
.I0(a[21]),
.I1(b[24]),
.I2(a[20]),
.I3(b[25]),
.I4(p_s0_o42_2),
.I5(1'b1));

wire p_s1_o43_2;
wire p_s1_o42_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o42_t96_z0_v1 (
.O6(p_s1_o43_2),
.O5(p_s1_o42_7),
.I0(a[19]),
.I1(b[26]),
.I2(a[18]),
.I3(b[27]),
.I4(p_s0_o42_3),
.I5(1'b1));

wire p_s1_o43_3;
wire p_s1_o42_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o42_t96_z0_v2 (
.O6(p_s1_o43_3),
.O5(p_s1_o42_8),
.I0(a[17]),
.I1(b[28]),
.I2(a[16]),
.I3(b[29]),
.I4(p_s0_o42_4),
.I5(1'b1));

wire p_s1_o43_4;
wire p_s1_o42_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o42_t96_z0_v3 (
.O6(p_s1_o43_4),
.O5(p_s1_o42_9),
.I0(a[15]),
.I1(b[30]),
.I2(a[14]),
.I3(b[31]),
.I4(p_s0_o42_5),
.I5(1'b1));

/////////STEP1----ORDER43////////////

wire p_s1_o44_0;
wire p_s1_o43_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o43_t97_z0_v0 (
.O6(p_s1_o44_0),
.O5(p_s1_o43_5),
.I0(a[25]),
.I1(b[21]),
.I2(a[24]),
.I3(b[22]),
.I4(p_s0_o43_0),
.I5(1'b1));

wire p_s1_o44_1;
wire p_s1_o43_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o43_t97_z0_v1 (
.O6(p_s1_o44_1),
.O5(p_s1_o43_6),
.I0(a[23]),
.I1(b[23]),
.I2(a[22]),
.I3(b[24]),
.I4(p_s0_o43_1),
.I5(1'b1));

wire p_s1_o44_2;
wire p_s1_o43_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o43_t97_z0_v2 (
.O6(p_s1_o44_2),
.O5(p_s1_o43_7),
.I0(a[21]),
.I1(b[25]),
.I2(a[20]),
.I3(b[26]),
.I4(p_s0_o43_2),
.I5(1'b1));

wire p_s1_o44_3;
wire p_s1_o43_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o43_t97_z0_v3 (
.O6(p_s1_o44_3),
.O5(p_s1_o43_8),
.I0(a[19]),
.I1(b[27]),
.I2(a[18]),
.I3(b[28]),
.I4(p_s0_o43_3),
.I5(1'b1));

wire p_s1_o44_4;
wire p_s1_o43_9;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o43_t97_z0_v4 (
.O6(p_s1_o44_4),
.O5(p_s1_o43_9),
.I0(a[17]),
.I1(b[29]),
.I2(a[16]),
.I3(b[30]),
.I4(p_s0_o43_4),
.I5(1'b1));

/////////STEP1----ORDER44////////////

wire p_s1_o45_0;
wire p_s1_o44_5;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s1_o44_t59_z0_v0 (
.O6(p_s1_o45_0),
.O5(p_s1_o44_5),
.I0(a[22]),
.I1(b[25]),
.I2(p_s0_o44_0),
.I3(p_s0_o44_1),
.I4(1'b0),
.I5(1'b1));

wire p_s1_o45_1;
wire p_s1_o44_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o44_t98_z0_v0 (
.O6(p_s1_o45_1),
.O5(p_s1_o44_6),
.I0(a[21]),
.I1(b[26]),
.I2(a[20]),
.I3(b[27]),
.I4(p_s0_o44_2),
.I5(1'b1));

wire p_s1_o45_2;
wire p_s1_o44_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o44_t98_z0_v1 (
.O6(p_s1_o45_2),
.O5(p_s1_o44_7),
.I0(a[19]),
.I1(b[28]),
.I2(a[18]),
.I3(b[29]),
.I4(p_s0_o44_3),
.I5(1'b1));

wire p_s1_o45_3;
wire p_s1_o44_8;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o44_t98_z0_v2 (
.O6(p_s1_o45_3),
.O5(p_s1_o44_8),
.I0(a[17]),
.I1(b[30]),
.I2(a[16]),
.I3(b[31]),
.I4(p_s0_o44_4),
.I5(1'b1));

/////////STEP1----ORDER45////////////

wire p_s1_o46_0;
wire p_s1_o45_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o45_t99_z0_v0 (
.O6(p_s1_o46_0),
.O5(p_s1_o45_4),
.I0(a[28]),
.I1(b[20]),
.I2(a[27]),
.I3(b[21]),
.I4(p_s0_o45_0),
.I5(1'b1));

wire p_s1_o46_1;
wire p_s1_o45_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o45_t99_z0_v1 (
.O6(p_s1_o46_1),
.O5(p_s1_o45_5),
.I0(a[26]),
.I1(b[22]),
.I2(a[25]),
.I3(b[23]),
.I4(p_s0_o45_1),
.I5(1'b1));

wire p_s1_o46_2;
wire p_s1_o45_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o45_t99_z0_v2 (
.O6(p_s1_o46_2),
.O5(p_s1_o45_6),
.I0(a[24]),
.I1(b[24]),
.I2(a[23]),
.I3(b[25]),
.I4(p_s0_o45_2),
.I5(1'b1));

wire p_s1_o46_3;
wire p_s1_o45_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o45_t99_z0_v3 (
.O6(p_s1_o46_3),
.O5(p_s1_o45_7),
.I0(a[22]),
.I1(b[26]),
.I2(a[21]),
.I3(b[27]),
.I4(p_s0_o45_3),
.I5(1'b1));

/////////STEP1----ORDER46////////////

wire p_s1_o47_0;
wire p_s1_o46_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o46_t100_z0_v0 (
.O6(p_s1_o47_0),
.O5(p_s1_o46_4),
.I0(a[25]),
.I1(b[24]),
.I2(a[24]),
.I3(b[25]),
.I4(p_s0_o46_0),
.I5(1'b1));

wire p_s1_o47_1;
wire p_s1_o46_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o46_t100_z0_v1 (
.O6(p_s1_o47_1),
.O5(p_s1_o46_5),
.I0(a[23]),
.I1(b[26]),
.I2(a[22]),
.I3(b[27]),
.I4(p_s0_o46_1),
.I5(1'b1));

wire p_s1_o47_2;
wire p_s1_o46_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o46_t100_z0_v2 (
.O6(p_s1_o47_2),
.O5(p_s1_o46_6),
.I0(a[21]),
.I1(b[28]),
.I2(a[20]),
.I3(b[29]),
.I4(p_s0_o46_2),
.I5(1'b1));

/////////STEP1----ORDER47////////////

wire p_s1_o48_0;
wire p_s1_o47_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o47_t101_z0_v0 (
.O6(p_s1_o48_0),
.O5(p_s1_o47_3),
.I0(a[28]),
.I1(b[22]),
.I2(a[27]),
.I3(b[23]),
.I4(p_s0_o47_0),
.I5(1'b1));

wire p_s1_o48_1;
wire p_s1_o47_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o47_t101_z0_v1 (
.O6(p_s1_o48_1),
.O5(p_s1_o47_4),
.I0(a[26]),
.I1(b[24]),
.I2(a[25]),
.I3(b[25]),
.I4(p_s0_o47_1),
.I5(1'b1));

wire p_s1_o48_2;
wire p_s1_o47_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o47_t101_z0_v2 (
.O6(p_s1_o48_2),
.O5(p_s1_o47_5),
.I0(a[24]),
.I1(b[26]),
.I2(a[23]),
.I3(b[27]),
.I4(p_s0_o47_2),
.I5(1'b1));

/////////STEP1----ORDER48////////////

wire p_s1_o49_0;
wire p_s1_o48_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o48_t102_z0_v0 (
.O6(p_s1_o49_0),
.O5(p_s1_o48_3),
.I0(a[25]),
.I1(b[26]),
.I2(a[24]),
.I3(b[27]),
.I4(p_s0_o48_0),
.I5(1'b1));

wire p_s1_o49_1;
wire p_s1_o48_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o48_t102_z0_v1 (
.O6(p_s1_o49_1),
.O5(p_s1_o48_4),
.I0(a[23]),
.I1(b[28]),
.I2(a[22]),
.I3(b[29]),
.I4(p_s0_o48_1),
.I5(1'b1));

wire p_s1_o49_2;
wire p_s1_o48_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o48_t102_z0_v2 (
.O6(p_s1_o49_2),
.O5(p_s1_o48_5),
.I0(a[21]),
.I1(b[30]),
.I2(a[20]),
.I3(b[31]),
.I4(p_s0_o48_2),
.I5(1'b1));

/////////STEP1----ORDER49////////////

wire p_s1_o50_0;
wire p_s1_o49_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o49_t103_z0_v0 (
.O6(p_s1_o50_0),
.O5(p_s1_o49_3),
.I0(a[31]),
.I1(b[21]),
.I2(a[30]),
.I3(b[22]),
.I4(p_s0_o49_0),
.I5(1'b1));

wire p_s1_o50_1;
wire p_s1_o49_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o49_t103_z0_v1 (
.O6(p_s1_o50_1),
.O5(p_s1_o49_4),
.I0(a[29]),
.I1(b[23]),
.I2(a[28]),
.I3(b[24]),
.I4(p_s0_o49_1),
.I5(1'b1));

/////////STEP1----ORDER50////////////

/////////STEP1----ORDER51////////////

wire p_s1_o52_0;
wire p_s1_o51_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o51_t104_z0_v0 (
.O6(p_s1_o52_0),
.O5(p_s1_o51_0),
.I0(a[28]),
.I1(b[26]),
.I2(a[27]),
.I3(b[27]),
.I4(p_s0_o51_0),
.I5(1'b1));

wire p_s1_o52_1;
wire p_s1_o51_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o51_t104_z0_v1 (
.O6(p_s1_o52_1),
.O5(p_s1_o51_1),
.I0(a[26]),
.I1(b[28]),
.I2(a[25]),
.I3(b[29]),
.I4(p_s0_o51_1),
.I5(1'b1));

/////////STEP1----ORDER52////////////

wire p_s1_o53_0;
wire p_s1_o52_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o52_t105_z0_v0 (
.O6(p_s1_o53_0),
.O5(p_s1_o52_2),
.I0(a[31]),
.I1(b[24]),
.I2(a[30]),
.I3(b[25]),
.I4(p_s0_o52_0),
.I5(1'b1));

/////////STEP1----ORDER53////////////

/////////STEP1----ORDER54////////////

wire p_s1_o55_0;
wire p_s1_o54_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o54_t106_z0_v0 (
.O6(p_s1_o55_0),
.O5(p_s1_o54_0),
.I0(a[28]),
.I1(b[29]),
.I2(a[27]),
.I3(b[30]),
.I4(p_s0_o54_0),
.I5(1'b1));

/////////STEP1----ORDER55////////////

wire p_s1_o56_0;
wire p_s1_o55_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o55_t107_z0_v0 (
.O6(p_s1_o56_0),
.O5(p_s1_o55_1),
.I0(a[31]),
.I1(b[27]),
.I2(a[30]),
.I3(b[28]),
.I4(p_s0_o55_0),
.I5(1'b1));

/////////STEP1----ORDER56////////////

/////////STEP1----ORDER57////////////

/////////STEP1----ORDER58////////////

/////////STEP1----ORDER59////////////

/////////STEP2----ORDER0////////////

/////////STEP2----ORDER1////////////

wire p_s2_o2_0;
wire p_s2_o1_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o1_t135_z0_v0 (
.O6(p_s2_o2_0),
.O5(p_s2_o1_0),
.I0(a[2]),
.I1(b[2]),
.I2(a[1]),
.I3(b[3]),
.I4(p_s1_o1_0),
.I5(1'b1));

/////////STEP2----ORDER2////////////

wire p_s2_o3_0;
wire p_s2_o2_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o2_t136_z0_v0 (
.O6(p_s2_o3_0),
.O5(p_s2_o2_1),
.I0(a[5]),
.I1(b[0]),
.I2(a[4]),
.I3(b[1]),
.I4(p_s1_o2_0),
.I5(1'b1));

/////////STEP2----ORDER3////////////

wire p_s2_o4_0;
wire p_s2_o3_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o3_t137_z0_v0 (
.O6(p_s2_o4_0),
.O5(p_s2_o3_1),
.I0(a[1]),
.I1(b[5]),
.I2(a[0]),
.I3(b[6]),
.I4(p_s1_o3_0),
.I5(1'b1));

/////////STEP2----ORDER4////////////

/////////STEP2----ORDER5////////////

wire p_s2_o6_0;
wire p_s2_o5_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o5_t138_z0_v0 (
.O6(p_s2_o6_0),
.O5(p_s2_o5_0),
.I0(a[6]),
.I1(b[2]),
.I2(a[5]),
.I3(b[3]),
.I4(p_s1_o5_0),
.I5(1'b1));

wire p_s2_o6_1;
wire p_s2_o5_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o5_t138_z0_v1 (
.O6(p_s2_o6_1),
.O5(p_s2_o5_1),
.I0(a[4]),
.I1(b[4]),
.I2(a[3]),
.I3(b[5]),
.I4(p_s1_o5_1),
.I5(1'b1));

wire p_s2_o6_2;
wire p_s2_o5_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o5_t138_z0_v2 (
.O6(p_s2_o6_2),
.O5(p_s2_o5_2),
.I0(a[2]),
.I1(b[6]),
.I2(a[1]),
.I3(b[7]),
.I4(p_s1_o5_2),
.I5(1'b1));

/////////STEP2----ORDER6////////////

wire p_s2_o7_0;
wire p_s2_o6_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o6_t139_z0_v0 (
.O6(p_s2_o7_0),
.O5(p_s2_o6_3),
.I0(a[9]),
.I1(b[0]),
.I2(a[8]),
.I3(b[1]),
.I4(p_s1_o6_0),
.I5(1'b1));

/////////STEP2----ORDER7////////////

wire p_s2_o8_0;
wire p_s2_o7_1;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o7_t130_z0_v0 (
.O6(p_s2_o8_0),
.O5(p_s2_o7_1),
.I0(a[0]),
.I1(b[10]),
.I2(p_s1_o7_0),
.I3(p_s1_o7_1),
.I4(1'b0),
.I5(1'b1));

/////////STEP2----ORDER8////////////

wire p_s2_o9_0;
wire p_s2_o8_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o8_t140_z0_v0 (
.O6(p_s2_o9_0),
.O5(p_s2_o8_1),
.I0(a[7]),
.I1(b[4]),
.I2(a[6]),
.I3(b[5]),
.I4(p_s1_o8_0),
.I5(1'b1));

wire p_s2_o9_1;
wire p_s2_o8_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o8_t140_z0_v1 (
.O6(p_s2_o9_1),
.O5(p_s2_o8_2),
.I0(a[5]),
.I1(b[6]),
.I2(a[4]),
.I3(b[7]),
.I4(p_s1_o8_1),
.I5(1'b1));

wire p_s2_o9_2;
wire p_s2_o8_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o8_t140_z0_v2 (
.O6(p_s2_o9_2),
.O5(p_s2_o8_3),
.I0(a[3]),
.I1(b[8]),
.I2(a[2]),
.I3(b[9]),
.I4(p_s1_o8_2),
.I5(1'b1));

wire p_s2_o9_3;
wire p_s2_o8_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o8_t140_z0_v3 (
.O6(p_s2_o9_3),
.O5(p_s2_o8_4),
.I0(a[1]),
.I1(b[10]),
.I2(a[0]),
.I3(b[11]),
.I4(p_s1_o8_3),
.I5(1'b1));

/////////STEP2----ORDER9////////////

wire p_s2_o10_0;
wire p_s2_o9_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o9_t141_z0_v0 (
.O6(p_s2_o10_0),
.O5(p_s2_o9_4),
.I0(a[7]),
.I1(b[5]),
.I2(a[6]),
.I3(b[6]),
.I4(p_s1_o9_0),
.I5(1'b1));

wire p_s2_o10_1;
wire p_s2_o9_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o9_t141_z0_v1 (
.O6(p_s2_o10_1),
.O5(p_s2_o9_5),
.I0(a[5]),
.I1(b[7]),
.I2(a[4]),
.I3(b[8]),
.I4(p_s1_o9_1),
.I5(1'b1));

wire p_s2_o10_2;
wire p_s2_o9_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o9_t141_z0_v2 (
.O6(p_s2_o10_2),
.O5(p_s2_o9_6),
.I0(a[3]),
.I1(b[9]),
.I2(a[2]),
.I3(b[10]),
.I4(p_s1_o9_2),
.I5(1'b1));

/////////STEP2----ORDER10////////////

wire p_s2_o11_0;
wire p_s2_o10_3;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s2_o10_t126_z0_v0 (
.O6(p_s2_o11_0),
.O5(p_s2_o10_3),
.I0(p_s1_o10_0),
.I1(p_s1_o10_1),
.I2(p_s1_o10_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o11_1;
wire p_s2_o10_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o10_t142_z0_v0 (
.O6(p_s2_o11_1),
.O5(p_s2_o10_4),
.I0(a[1]),
.I1(b[12]),
.I2(a[0]),
.I3(b[13]),
.I4(p_s1_o10_3),
.I5(1'b1));

/////////STEP2----ORDER11////////////

wire p_s2_o12_0;
wire p_s2_o11_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o11_t143_z0_v0 (
.O6(p_s2_o12_0),
.O5(p_s2_o11_2),
.I0(a[1]),
.I1(b[13]),
.I2(a[0]),
.I3(b[14]),
.I4(p_s1_o11_0),
.I5(1'b1));

wire p_s2_o11_3;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o11_t155_z0_v0 (
.O6(p_s2_o11_3),
.O5(),
.I0(p_s1_o11_1),
.I1(p_s1_o11_2),
.I2(p_s1_o11_3),
.I3(p_s1_o11_4),
.I4(p_s1_o11_5),
.I5(p_s1_o11_6));

wire p_s2_o12_1;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o11_t155_z1_v0 (
.O6(p_s2_o12_1),
.O5(),
.I0(p_s1_o11_1),
.I1(p_s1_o11_2),
.I2(p_s1_o11_3),
.I3(p_s1_o11_4),
.I4(p_s1_o11_5),
.I5(p_s1_o11_6));

wire p_s2_o13_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o11_t155_z2_v0 (
.O6(p_s2_o13_0),
.O5(),
.I0(p_s1_o11_1),
.I1(p_s1_o11_2),
.I2(p_s1_o11_3),
.I3(p_s1_o11_4),
.I4(p_s1_o11_5),
.I5(p_s1_o11_6));

/////////STEP2----ORDER12////////////

wire p_s2_o13_1;
wire p_s2_o12_2;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o12_t131_z0_v0 (
.O6(p_s2_o13_1),
.O5(p_s2_o12_2),
.I0(a[7]),
.I1(b[8]),
.I2(p_s1_o12_0),
.I3(p_s1_o12_1),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o13_2;
wire p_s2_o12_3;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o12_t131_z0_v1 (
.O6(p_s2_o13_2),
.O5(p_s2_o12_3),
.I0(a[6]),
.I1(b[9]),
.I2(p_s1_o12_2),
.I3(p_s1_o12_3),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o13_3;
wire p_s2_o12_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o12_t144_z0_v0 (
.O6(p_s2_o13_3),
.O5(p_s2_o12_4),
.I0(a[5]),
.I1(b[10]),
.I2(a[4]),
.I3(b[11]),
.I4(p_s1_o12_4),
.I5(1'b1));

wire p_s2_o13_4;
wire p_s2_o12_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o12_t144_z0_v1 (
.O6(p_s2_o13_4),
.O5(p_s2_o12_5),
.I0(a[3]),
.I1(b[12]),
.I2(a[2]),
.I3(b[13]),
.I4(p_s1_o12_5),
.I5(1'b1));

wire p_s2_o13_5;
wire p_s2_o12_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o12_t144_z0_v2 (
.O6(p_s2_o13_5),
.O5(p_s2_o12_6),
.I0(a[1]),
.I1(b[14]),
.I2(a[0]),
.I3(b[15]),
.I4(p_s1_o12_6),
.I5(1'b1));

/////////STEP2----ORDER13////////////

wire p_s2_o13_6;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o13_t167_z0_v0 (
.O6(p_s2_o13_6),
.O5(),
.I0(p_s1_o13_0),
.I1(p_s1_o13_1),
.I2(p_s1_o13_2),
.I3(p_s1_o13_3),
.I4(p_s1_o13_4),
.I5(p_s1_o14_0));

wire p_s2_o14_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o13_t167_z1_v0 (
.O6(p_s2_o14_0),
.O5(),
.I0(p_s1_o13_0),
.I1(p_s1_o13_1),
.I2(p_s1_o13_2),
.I3(p_s1_o13_3),
.I4(p_s1_o13_4),
.I5(p_s1_o14_0));

wire p_s2_o15_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o13_t167_z2_v0 (
.O6(p_s2_o15_0),
.O5(),
.I0(p_s1_o13_0),
.I1(p_s1_o13_1),
.I2(p_s1_o13_2),
.I3(p_s1_o13_3),
.I4(p_s1_o13_4),
.I5(p_s1_o14_0));

/////////STEP2----ORDER14////////////

wire p_s2_o14_1;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o14_t156_z0_v0 (
.O6(p_s2_o14_1),
.O5(),
.I0(p_s1_o14_1),
.I1(p_s1_o14_2),
.I2(p_s1_o14_3),
.I3(p_s1_o14_4),
.I4(p_s1_o14_5),
.I5(p_s1_o14_6));

wire p_s2_o15_1;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o14_t156_z1_v0 (
.O6(p_s2_o15_1),
.O5(),
.I0(p_s1_o14_1),
.I1(p_s1_o14_2),
.I2(p_s1_o14_3),
.I3(p_s1_o14_4),
.I4(p_s1_o14_5),
.I5(p_s1_o14_6));

wire p_s2_o16_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o14_t156_z2_v0 (
.O6(p_s2_o16_0),
.O5(),
.I0(p_s1_o14_1),
.I1(p_s1_o14_2),
.I2(p_s1_o14_3),
.I3(p_s1_o14_4),
.I4(p_s1_o14_5),
.I5(p_s1_o14_6));

/////////STEP2----ORDER15////////////

wire p_s2_o15_2;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o15_t157_z0_v0 (
.O6(p_s2_o15_2),
.O5(),
.I0(p_s1_o15_0),
.I1(p_s1_o15_1),
.I2(p_s1_o15_2),
.I3(p_s1_o15_3),
.I4(p_s1_o15_4),
.I5(p_s1_o15_5));

wire p_s2_o16_1;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o15_t157_z1_v0 (
.O6(p_s2_o16_1),
.O5(),
.I0(p_s1_o15_0),
.I1(p_s1_o15_1),
.I2(p_s1_o15_2),
.I3(p_s1_o15_3),
.I4(p_s1_o15_4),
.I5(p_s1_o15_5));

wire p_s2_o17_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o15_t157_z2_v0 (
.O6(p_s2_o17_0),
.O5(),
.I0(p_s1_o15_0),
.I1(p_s1_o15_1),
.I2(p_s1_o15_2),
.I3(p_s1_o15_3),
.I4(p_s1_o15_4),
.I5(p_s1_o15_5));

wire p_s2_o15_3;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o15_t157_z0_v1 (
.O6(p_s2_o15_3),
.O5(),
.I0(p_s1_o15_6),
.I1(p_s1_o15_7),
.I2(p_s1_o15_8),
.I3(p_s1_o15_9),
.I4(p_s1_o15_10),
.I5(p_s1_o15_11));

wire p_s2_o16_2;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o15_t157_z1_v1 (
.O6(p_s2_o16_2),
.O5(),
.I0(p_s1_o15_6),
.I1(p_s1_o15_7),
.I2(p_s1_o15_8),
.I3(p_s1_o15_9),
.I4(p_s1_o15_10),
.I5(p_s1_o15_11));

wire p_s2_o17_1;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o15_t157_z2_v1 (
.O6(p_s2_o17_1),
.O5(),
.I0(p_s1_o15_6),
.I1(p_s1_o15_7),
.I2(p_s1_o15_8),
.I3(p_s1_o15_9),
.I4(p_s1_o15_10),
.I5(p_s1_o15_11));

/////////STEP2----ORDER16////////////

wire p_s2_o17_2;
wire p_s2_o16_3;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s2_o16_t127_z0_v0 (
.O6(p_s2_o17_2),
.O5(p_s2_o16_3),
.I0(p_s1_o16_0),
.I1(p_s1_o16_1),
.I2(p_s1_o16_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o17_3;
wire p_s2_o16_4;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o16_t132_z0_v0 (
.O6(p_s2_o17_3),
.O5(p_s2_o16_4),
.I0(a[0]),
.I1(b[19]),
.I2(p_s1_o16_3),
.I3(p_s1_o16_4),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o16_5;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o16_t158_z0_v0 (
.O6(p_s2_o16_5),
.O5(),
.I0(p_s1_o16_5),
.I1(p_s1_o16_6),
.I2(p_s1_o16_7),
.I3(p_s1_o16_8),
.I4(p_s1_o16_9),
.I5(p_s0_o16_5));

wire p_s2_o17_4;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o16_t158_z1_v0 (
.O6(p_s2_o17_4),
.O5(),
.I0(p_s1_o16_5),
.I1(p_s1_o16_6),
.I2(p_s1_o16_7),
.I3(p_s1_o16_8),
.I4(p_s1_o16_9),
.I5(p_s0_o16_5));

wire p_s2_o18_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o16_t158_z2_v0 (
.O6(p_s2_o18_0),
.O5(),
.I0(p_s1_o16_5),
.I1(p_s1_o16_6),
.I2(p_s1_o16_7),
.I3(p_s1_o16_8),
.I4(p_s1_o16_9),
.I5(p_s0_o16_5));

/////////STEP2----ORDER17////////////

wire p_s2_o17_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o17_t168_z0_v0 (
.O6(p_s2_o17_5),
.O5(),
.I0(p_s1_o17_0),
.I1(p_s1_o17_1),
.I2(p_s1_o17_2),
.I3(p_s1_o17_3),
.I4(p_s1_o17_4),
.I5(p_s1_o18_0));

wire p_s2_o18_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o17_t168_z1_v0 (
.O6(p_s2_o18_1),
.O5(),
.I0(p_s1_o17_0),
.I1(p_s1_o17_1),
.I2(p_s1_o17_2),
.I3(p_s1_o17_3),
.I4(p_s1_o17_4),
.I5(p_s1_o18_0));

wire p_s2_o19_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o17_t168_z2_v0 (
.O6(p_s2_o19_0),
.O5(),
.I0(p_s1_o17_0),
.I1(p_s1_o17_1),
.I2(p_s1_o17_2),
.I3(p_s1_o17_3),
.I4(p_s1_o17_4),
.I5(p_s1_o18_0));

wire p_s2_o17_6;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o17_t168_z0_v1 (
.O6(p_s2_o17_6),
.O5(),
.I0(p_s1_o17_5),
.I1(p_s1_o17_6),
.I2(p_s1_o17_7),
.I3(p_s1_o17_8),
.I4(p_s1_o17_9),
.I5(p_s1_o18_1));

wire p_s2_o18_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o17_t168_z1_v1 (
.O6(p_s2_o18_2),
.O5(),
.I0(p_s1_o17_5),
.I1(p_s1_o17_6),
.I2(p_s1_o17_7),
.I3(p_s1_o17_8),
.I4(p_s1_o17_9),
.I5(p_s1_o18_1));

wire p_s2_o19_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o17_t168_z2_v1 (
.O6(p_s2_o19_1),
.O5(),
.I0(p_s1_o17_5),
.I1(p_s1_o17_6),
.I2(p_s1_o17_7),
.I3(p_s1_o17_8),
.I4(p_s1_o17_9),
.I5(p_s1_o18_1));

/////////STEP2----ORDER18////////////

wire p_s2_o18_3;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o18_t159_z0_v0 (
.O6(p_s2_o18_3),
.O5(),
.I0(p_s1_o18_2),
.I1(p_s1_o18_3),
.I2(p_s1_o18_4),
.I3(p_s1_o18_5),
.I4(p_s1_o18_6),
.I5(p_s1_o18_7));

wire p_s2_o19_2;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o18_t159_z1_v0 (
.O6(p_s2_o19_2),
.O5(),
.I0(p_s1_o18_2),
.I1(p_s1_o18_3),
.I2(p_s1_o18_4),
.I3(p_s1_o18_5),
.I4(p_s1_o18_6),
.I5(p_s1_o18_7));

wire p_s2_o20_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o18_t159_z2_v0 (
.O6(p_s2_o20_0),
.O5(),
.I0(p_s1_o18_2),
.I1(p_s1_o18_3),
.I2(p_s1_o18_4),
.I3(p_s1_o18_5),
.I4(p_s1_o18_6),
.I5(p_s1_o18_7));

wire p_s2_o18_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o18_t169_z0_v0 (
.O6(p_s2_o18_4),
.O5(),
.I0(p_s1_o18_8),
.I1(p_s1_o18_9),
.I2(p_s1_o18_10),
.I3(p_s0_o18_5),
.I4(p_s0_o18_6),
.I5(p_s1_o19_0));

wire p_s2_o19_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o18_t169_z1_v0 (
.O6(p_s2_o19_3),
.O5(),
.I0(p_s1_o18_8),
.I1(p_s1_o18_9),
.I2(p_s1_o18_10),
.I3(p_s0_o18_5),
.I4(p_s0_o18_6),
.I5(p_s1_o19_0));

wire p_s2_o20_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o18_t169_z2_v0 (
.O6(p_s2_o20_1),
.O5(),
.I0(p_s1_o18_8),
.I1(p_s1_o18_9),
.I2(p_s1_o18_10),
.I3(p_s0_o18_5),
.I4(p_s0_o18_6),
.I5(p_s1_o19_0));

/////////STEP2----ORDER19////////////

wire p_s2_o19_4;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o19_t160_z0_v0 (
.O6(p_s2_o19_4),
.O5(),
.I0(p_s1_o19_1),
.I1(p_s1_o19_2),
.I2(p_s1_o19_3),
.I3(p_s1_o19_4),
.I4(p_s1_o19_5),
.I5(p_s1_o19_6));

wire p_s2_o20_2;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o19_t160_z1_v0 (
.O6(p_s2_o20_2),
.O5(),
.I0(p_s1_o19_1),
.I1(p_s1_o19_2),
.I2(p_s1_o19_3),
.I3(p_s1_o19_4),
.I4(p_s1_o19_5),
.I5(p_s1_o19_6));

wire p_s2_o21_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o19_t160_z2_v0 (
.O6(p_s2_o21_0),
.O5(),
.I0(p_s1_o19_1),
.I1(p_s1_o19_2),
.I2(p_s1_o19_3),
.I3(p_s1_o19_4),
.I4(p_s1_o19_5),
.I5(p_s1_o19_6));

wire p_s2_o19_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o19_t170_z0_v0 (
.O6(p_s2_o19_5),
.O5(),
.I0(p_s1_o19_7),
.I1(p_s1_o19_8),
.I2(p_s1_o19_9),
.I3(p_s1_o19_10),
.I4(p_s1_o19_11),
.I5(p_s1_o20_0));

wire p_s2_o20_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o19_t170_z1_v0 (
.O6(p_s2_o20_3),
.O5(),
.I0(p_s1_o19_7),
.I1(p_s1_o19_8),
.I2(p_s1_o19_9),
.I3(p_s1_o19_10),
.I4(p_s1_o19_11),
.I5(p_s1_o20_0));

wire p_s2_o21_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o19_t170_z2_v0 (
.O6(p_s2_o21_1),
.O5(),
.I0(p_s1_o19_7),
.I1(p_s1_o19_8),
.I2(p_s1_o19_9),
.I3(p_s1_o19_10),
.I4(p_s1_o19_11),
.I5(p_s1_o20_0));

/////////STEP2----ORDER20////////////

wire p_s2_o20_4;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o20_t161_z0_v0 (
.O6(p_s2_o20_4),
.O5(),
.I0(p_s1_o20_1),
.I1(p_s1_o20_2),
.I2(p_s1_o20_3),
.I3(p_s1_o20_4),
.I4(p_s1_o20_5),
.I5(p_s1_o20_6));

wire p_s2_o21_2;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o20_t161_z1_v0 (
.O6(p_s2_o21_2),
.O5(),
.I0(p_s1_o20_1),
.I1(p_s1_o20_2),
.I2(p_s1_o20_3),
.I3(p_s1_o20_4),
.I4(p_s1_o20_5),
.I5(p_s1_o20_6));

wire p_s2_o22_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o20_t161_z2_v0 (
.O6(p_s2_o22_0),
.O5(),
.I0(p_s1_o20_1),
.I1(p_s1_o20_2),
.I2(p_s1_o20_3),
.I3(p_s1_o20_4),
.I4(p_s1_o20_5),
.I5(p_s1_o20_6));

wire p_s2_o20_5;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o20_t161_z0_v1 (
.O6(p_s2_o20_5),
.O5(),
.I0(p_s1_o20_7),
.I1(p_s1_o20_8),
.I2(p_s1_o20_9),
.I3(p_s1_o20_10),
.I4(p_s0_o20_7),
.I5(p_s0_o20_8));

wire p_s2_o21_3;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o20_t161_z1_v1 (
.O6(p_s2_o21_3),
.O5(),
.I0(p_s1_o20_7),
.I1(p_s1_o20_8),
.I2(p_s1_o20_9),
.I3(p_s1_o20_10),
.I4(p_s0_o20_7),
.I5(p_s0_o20_8));

wire p_s2_o22_1;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o20_t161_z2_v1 (
.O6(p_s2_o22_1),
.O5(),
.I0(p_s1_o20_7),
.I1(p_s1_o20_8),
.I2(p_s1_o20_9),
.I3(p_s1_o20_10),
.I4(p_s0_o20_7),
.I5(p_s0_o20_8));

/////////STEP2----ORDER21////////////

wire p_s2_o21_4;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o21_t162_z0_v0 (
.O6(p_s2_o21_4),
.O5(),
.I0(p_s1_o21_0),
.I1(p_s1_o21_1),
.I2(p_s1_o21_2),
.I3(p_s1_o21_3),
.I4(p_s1_o21_4),
.I5(p_s1_o21_5));

wire p_s2_o22_2;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o21_t162_z1_v0 (
.O6(p_s2_o22_2),
.O5(),
.I0(p_s1_o21_0),
.I1(p_s1_o21_1),
.I2(p_s1_o21_2),
.I3(p_s1_o21_3),
.I4(p_s1_o21_4),
.I5(p_s1_o21_5));

wire p_s2_o23_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o21_t162_z2_v0 (
.O6(p_s2_o23_0),
.O5(),
.I0(p_s1_o21_0),
.I1(p_s1_o21_1),
.I2(p_s1_o21_2),
.I3(p_s1_o21_3),
.I4(p_s1_o21_4),
.I5(p_s1_o21_5));

wire p_s2_o21_5;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o21_t162_z0_v1 (
.O6(p_s2_o21_5),
.O5(),
.I0(p_s1_o21_6),
.I1(p_s1_o21_7),
.I2(p_s1_o21_8),
.I3(p_s1_o21_9),
.I4(p_s1_o21_10),
.I5(p_s1_o21_11));

wire p_s2_o22_3;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o21_t162_z1_v1 (
.O6(p_s2_o22_3),
.O5(),
.I0(p_s1_o21_6),
.I1(p_s1_o21_7),
.I2(p_s1_o21_8),
.I3(p_s1_o21_9),
.I4(p_s1_o21_10),
.I5(p_s1_o21_11));

wire p_s2_o23_1;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o21_t162_z2_v1 (
.O6(p_s2_o23_1),
.O5(),
.I0(p_s1_o21_6),
.I1(p_s1_o21_7),
.I2(p_s1_o21_8),
.I3(p_s1_o21_9),
.I4(p_s1_o21_10),
.I5(p_s1_o21_11));

/////////STEP2----ORDER22////////////

wire p_s2_o22_4;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o22_t163_z0_v0 (
.O6(p_s2_o22_4),
.O5(),
.I0(p_s1_o22_0),
.I1(p_s1_o22_1),
.I2(p_s1_o22_2),
.I3(p_s1_o22_3),
.I4(p_s1_o22_4),
.I5(p_s1_o22_5));

wire p_s2_o23_2;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o22_t163_z1_v0 (
.O6(p_s2_o23_2),
.O5(),
.I0(p_s1_o22_0),
.I1(p_s1_o22_1),
.I2(p_s1_o22_2),
.I3(p_s1_o22_3),
.I4(p_s1_o22_4),
.I5(p_s1_o22_5));

wire p_s2_o24_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o22_t163_z2_v0 (
.O6(p_s2_o24_0),
.O5(),
.I0(p_s1_o22_0),
.I1(p_s1_o22_1),
.I2(p_s1_o22_2),
.I3(p_s1_o22_3),
.I4(p_s1_o22_4),
.I5(p_s1_o22_5));

wire p_s2_o22_5;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o22_t163_z0_v1 (
.O6(p_s2_o22_5),
.O5(),
.I0(p_s1_o22_6),
.I1(p_s1_o22_7),
.I2(p_s1_o22_8),
.I3(p_s1_o22_9),
.I4(p_s1_o22_10),
.I5(p_s1_o22_11));

wire p_s2_o23_3;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o22_t163_z1_v1 (
.O6(p_s2_o23_3),
.O5(),
.I0(p_s1_o22_6),
.I1(p_s1_o22_7),
.I2(p_s1_o22_8),
.I3(p_s1_o22_9),
.I4(p_s1_o22_10),
.I5(p_s1_o22_11));

wire p_s2_o24_1;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o22_t163_z2_v1 (
.O6(p_s2_o24_1),
.O5(),
.I0(p_s1_o22_6),
.I1(p_s1_o22_7),
.I2(p_s1_o22_8),
.I3(p_s1_o22_9),
.I4(p_s1_o22_10),
.I5(p_s1_o22_11));

/////////STEP2----ORDER23////////////

wire p_s2_o23_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o23_t171_z0_v0 (
.O6(p_s2_o23_4),
.O5(),
.I0(p_s1_o23_0),
.I1(p_s1_o23_1),
.I2(p_s1_o23_2),
.I3(p_s1_o23_3),
.I4(p_s1_o23_4),
.I5(p_s1_o24_0));

wire p_s2_o24_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o23_t171_z1_v0 (
.O6(p_s2_o24_2),
.O5(),
.I0(p_s1_o23_0),
.I1(p_s1_o23_1),
.I2(p_s1_o23_2),
.I3(p_s1_o23_3),
.I4(p_s1_o23_4),
.I5(p_s1_o24_0));

wire p_s2_o25_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o23_t171_z2_v0 (
.O6(p_s2_o25_0),
.O5(),
.I0(p_s1_o23_0),
.I1(p_s1_o23_1),
.I2(p_s1_o23_2),
.I3(p_s1_o23_3),
.I4(p_s1_o23_4),
.I5(p_s1_o24_0));

wire p_s2_o23_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o23_t171_z0_v1 (
.O6(p_s2_o23_5),
.O5(),
.I0(p_s1_o23_5),
.I1(p_s1_o23_6),
.I2(p_s1_o23_7),
.I3(p_s1_o23_8),
.I4(p_s1_o23_9),
.I5(p_s1_o24_1));

wire p_s2_o24_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o23_t171_z1_v1 (
.O6(p_s2_o24_3),
.O5(),
.I0(p_s1_o23_5),
.I1(p_s1_o23_6),
.I2(p_s1_o23_7),
.I3(p_s1_o23_8),
.I4(p_s1_o23_9),
.I5(p_s1_o24_1));

wire p_s2_o25_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o23_t171_z2_v1 (
.O6(p_s2_o25_1),
.O5(),
.I0(p_s1_o23_5),
.I1(p_s1_o23_6),
.I2(p_s1_o23_7),
.I3(p_s1_o23_8),
.I4(p_s1_o23_9),
.I5(p_s1_o24_1));

/////////STEP2----ORDER24////////////

wire p_s2_o24_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o24_t172_z0_v0 (
.O6(p_s2_o24_4),
.O5(),
.I0(p_s1_o24_2),
.I1(p_s1_o24_3),
.I2(p_s1_o24_4),
.I3(p_s1_o24_5),
.I4(p_s1_o24_6),
.I5(p_s1_o25_0));

wire p_s2_o25_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o24_t172_z1_v0 (
.O6(p_s2_o25_2),
.O5(),
.I0(p_s1_o24_2),
.I1(p_s1_o24_3),
.I2(p_s1_o24_4),
.I3(p_s1_o24_5),
.I4(p_s1_o24_6),
.I5(p_s1_o25_0));

wire p_s2_o26_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o24_t172_z2_v0 (
.O6(p_s2_o26_0),
.O5(),
.I0(p_s1_o24_2),
.I1(p_s1_o24_3),
.I2(p_s1_o24_4),
.I3(p_s1_o24_5),
.I4(p_s1_o24_6),
.I5(p_s1_o25_0));

wire p_s2_o24_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o24_t172_z0_v1 (
.O6(p_s2_o24_5),
.O5(),
.I0(p_s1_o24_7),
.I1(p_s1_o24_8),
.I2(p_s1_o24_9),
.I3(p_s1_o24_10),
.I4(p_s1_o24_11),
.I5(p_s1_o25_1));

wire p_s2_o25_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o24_t172_z1_v1 (
.O6(p_s2_o25_3),
.O5(),
.I0(p_s1_o24_7),
.I1(p_s1_o24_8),
.I2(p_s1_o24_9),
.I3(p_s1_o24_10),
.I4(p_s1_o24_11),
.I5(p_s1_o25_1));

wire p_s2_o26_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o24_t172_z2_v1 (
.O6(p_s2_o26_1),
.O5(),
.I0(p_s1_o24_7),
.I1(p_s1_o24_8),
.I2(p_s1_o24_9),
.I3(p_s1_o24_10),
.I4(p_s1_o24_11),
.I5(p_s1_o25_1));

/////////STEP2----ORDER25////////////

wire p_s2_o25_4;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o25_t164_z0_v0 (
.O6(p_s2_o25_4),
.O5(),
.I0(p_s1_o25_2),
.I1(p_s1_o25_3),
.I2(p_s1_o25_4),
.I3(p_s1_o25_5),
.I4(p_s1_o25_6),
.I5(p_s1_o25_7));

wire p_s2_o26_2;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o25_t164_z1_v0 (
.O6(p_s2_o26_2),
.O5(),
.I0(p_s1_o25_2),
.I1(p_s1_o25_3),
.I2(p_s1_o25_4),
.I3(p_s1_o25_5),
.I4(p_s1_o25_6),
.I5(p_s1_o25_7));

wire p_s2_o27_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o25_t164_z2_v0 (
.O6(p_s2_o27_0),
.O5(),
.I0(p_s1_o25_2),
.I1(p_s1_o25_3),
.I2(p_s1_o25_4),
.I3(p_s1_o25_5),
.I4(p_s1_o25_6),
.I5(p_s1_o25_7));

wire p_s2_o25_5;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o25_t164_z0_v1 (
.O6(p_s2_o25_5),
.O5(),
.I0(p_s1_o25_8),
.I1(p_s1_o25_9),
.I2(p_s1_o25_10),
.I3(p_s1_o25_11),
.I4(p_s1_o25_12),
.I5(p_s1_o25_13));

wire p_s2_o26_3;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o25_t164_z1_v1 (
.O6(p_s2_o26_3),
.O5(),
.I0(p_s1_o25_8),
.I1(p_s1_o25_9),
.I2(p_s1_o25_10),
.I3(p_s1_o25_11),
.I4(p_s1_o25_12),
.I5(p_s1_o25_13));

wire p_s2_o27_1;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o25_t164_z2_v1 (
.O6(p_s2_o27_1),
.O5(),
.I0(p_s1_o25_8),
.I1(p_s1_o25_9),
.I2(p_s1_o25_10),
.I3(p_s1_o25_11),
.I4(p_s1_o25_12),
.I5(p_s1_o25_13));

/////////STEP2----ORDER26////////////

wire p_s2_o26_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o26_t173_z0_v0 (
.O6(p_s2_o26_4),
.O5(),
.I0(p_s1_o26_0),
.I1(p_s1_o26_1),
.I2(p_s1_o26_2),
.I3(p_s1_o26_3),
.I4(p_s1_o26_4),
.I5(p_s1_o27_0));

wire p_s2_o27_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o26_t173_z1_v0 (
.O6(p_s2_o27_2),
.O5(),
.I0(p_s1_o26_0),
.I1(p_s1_o26_1),
.I2(p_s1_o26_2),
.I3(p_s1_o26_3),
.I4(p_s1_o26_4),
.I5(p_s1_o27_0));

wire p_s2_o28_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o26_t173_z2_v0 (
.O6(p_s2_o28_0),
.O5(),
.I0(p_s1_o26_0),
.I1(p_s1_o26_1),
.I2(p_s1_o26_2),
.I3(p_s1_o26_3),
.I4(p_s1_o26_4),
.I5(p_s1_o27_0));

wire p_s2_o26_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o26_t173_z0_v1 (
.O6(p_s2_o26_5),
.O5(),
.I0(p_s1_o26_5),
.I1(p_s1_o26_6),
.I2(p_s1_o26_7),
.I3(p_s1_o26_8),
.I4(p_s1_o26_9),
.I5(p_s1_o27_1));

wire p_s2_o27_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o26_t173_z1_v1 (
.O6(p_s2_o27_3),
.O5(),
.I0(p_s1_o26_5),
.I1(p_s1_o26_6),
.I2(p_s1_o26_7),
.I3(p_s1_o26_8),
.I4(p_s1_o26_9),
.I5(p_s1_o27_1));

wire p_s2_o28_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o26_t173_z2_v1 (
.O6(p_s2_o28_1),
.O5(),
.I0(p_s1_o26_5),
.I1(p_s1_o26_6),
.I2(p_s1_o26_7),
.I3(p_s1_o26_8),
.I4(p_s1_o26_9),
.I5(p_s1_o27_1));

wire p_s2_o26_6;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o26_t173_z0_v2 (
.O6(p_s2_o26_6),
.O5(),
.I0(p_s1_o26_10),
.I1(p_s1_o26_11),
.I2(p_s1_o26_12),
.I3(p_s1_o26_13),
.I4(p_s0_o26_12),
.I5(p_s1_o27_2));

wire p_s2_o27_4;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o26_t173_z1_v2 (
.O6(p_s2_o27_4),
.O5(),
.I0(p_s1_o26_10),
.I1(p_s1_o26_11),
.I2(p_s1_o26_12),
.I3(p_s1_o26_13),
.I4(p_s0_o26_12),
.I5(p_s1_o27_2));

wire p_s2_o28_2;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o26_t173_z2_v2 (
.O6(p_s2_o28_2),
.O5(),
.I0(p_s1_o26_10),
.I1(p_s1_o26_11),
.I2(p_s1_o26_12),
.I3(p_s1_o26_13),
.I4(p_s0_o26_12),
.I5(p_s1_o27_2));

/////////STEP2----ORDER27////////////

wire p_s2_o27_5;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o27_t165_z0_v0 (
.O6(p_s2_o27_5),
.O5(),
.I0(p_s1_o27_3),
.I1(p_s1_o27_4),
.I2(p_s1_o27_5),
.I3(p_s1_o27_6),
.I4(p_s0_o27_17),
.I5(p_s0_o27_18));

wire p_s2_o28_3;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o27_t165_z1_v0 (
.O6(p_s2_o28_3),
.O5(),
.I0(p_s1_o27_3),
.I1(p_s1_o27_4),
.I2(p_s1_o27_5),
.I3(p_s1_o27_6),
.I4(p_s0_o27_17),
.I5(p_s0_o27_18));

wire p_s2_o29_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o27_t165_z2_v0 (
.O6(p_s2_o29_0),
.O5(),
.I0(p_s1_o27_3),
.I1(p_s1_o27_4),
.I2(p_s1_o27_5),
.I3(p_s1_o27_6),
.I4(p_s0_o27_17),
.I5(p_s0_o27_18));

/////////STEP2----ORDER28////////////

wire p_s2_o28_4;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s2_o28_t166_z0_v0 (
.O6(p_s2_o28_4),
.O5(),
.I0(p_s1_o28_0),
.I1(p_s1_o28_1),
.I2(p_s1_o28_2),
.I3(p_s1_o28_3),
.I4(p_s1_o28_4),
.I5(p_s1_o28_5));

wire p_s2_o29_1;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s2_o28_t166_z1_v0 (
.O6(p_s2_o29_1),
.O5(),
.I0(p_s1_o28_0),
.I1(p_s1_o28_1),
.I2(p_s1_o28_2),
.I3(p_s1_o28_3),
.I4(p_s1_o28_4),
.I5(p_s1_o28_5));

wire p_s2_o30_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s2_o28_t166_z2_v0 (
.O6(p_s2_o30_0),
.O5(),
.I0(p_s1_o28_0),
.I1(p_s1_o28_1),
.I2(p_s1_o28_2),
.I3(p_s1_o28_3),
.I4(p_s1_o28_4),
.I5(p_s1_o28_5));

wire p_s2_o28_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o28_t174_z0_v0 (
.O6(p_s2_o28_5),
.O5(),
.I0(p_s1_o28_6),
.I1(p_s1_o28_7),
.I2(p_s1_o28_8),
.I3(p_s1_o28_9),
.I4(p_s1_o28_10),
.I5(p_s1_o29_0));

wire p_s2_o29_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o28_t174_z1_v0 (
.O6(p_s2_o29_2),
.O5(),
.I0(p_s1_o28_6),
.I1(p_s1_o28_7),
.I2(p_s1_o28_8),
.I3(p_s1_o28_9),
.I4(p_s1_o28_10),
.I5(p_s1_o29_0));

wire p_s2_o30_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o28_t174_z2_v0 (
.O6(p_s2_o30_1),
.O5(),
.I0(p_s1_o28_6),
.I1(p_s1_o28_7),
.I2(p_s1_o28_8),
.I3(p_s1_o28_9),
.I4(p_s1_o28_10),
.I5(p_s1_o29_0));

/////////STEP2----ORDER29////////////

wire p_s2_o29_3;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o29_t175_z0_v0 (
.O6(p_s2_o29_3),
.O5(),
.I0(p_s1_o29_1),
.I1(p_s1_o29_2),
.I2(p_s1_o29_3),
.I3(p_s1_o29_4),
.I4(p_s1_o29_5),
.I5(p_s1_o30_0));

wire p_s2_o30_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o29_t175_z1_v0 (
.O6(p_s2_o30_2),
.O5(),
.I0(p_s1_o29_1),
.I1(p_s1_o29_2),
.I2(p_s1_o29_3),
.I3(p_s1_o29_4),
.I4(p_s1_o29_5),
.I5(p_s1_o30_0));

wire p_s2_o31_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o29_t175_z2_v0 (
.O6(p_s2_o31_0),
.O5(),
.I0(p_s1_o29_1),
.I1(p_s1_o29_2),
.I2(p_s1_o29_3),
.I3(p_s1_o29_4),
.I4(p_s1_o29_5),
.I5(p_s1_o30_0));

wire p_s2_o29_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o29_t175_z0_v1 (
.O6(p_s2_o29_4),
.O5(),
.I0(p_s1_o29_6),
.I1(p_s1_o29_7),
.I2(p_s1_o29_8),
.I3(p_s1_o29_9),
.I4(p_s1_o29_10),
.I5(p_s1_o30_1));

wire p_s2_o30_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o29_t175_z1_v1 (
.O6(p_s2_o30_3),
.O5(),
.I0(p_s1_o29_6),
.I1(p_s1_o29_7),
.I2(p_s1_o29_8),
.I3(p_s1_o29_9),
.I4(p_s1_o29_10),
.I5(p_s1_o30_1));

wire p_s2_o31_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o29_t175_z2_v1 (
.O6(p_s2_o31_1),
.O5(),
.I0(p_s1_o29_6),
.I1(p_s1_o29_7),
.I2(p_s1_o29_8),
.I3(p_s1_o29_9),
.I4(p_s1_o29_10),
.I5(p_s1_o30_1));

/////////STEP2----ORDER30////////////

wire p_s2_o30_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o30_t176_z0_v0 (
.O6(p_s2_o30_4),
.O5(),
.I0(p_s1_o30_2),
.I1(p_s1_o30_3),
.I2(p_s1_o30_4),
.I3(p_s1_o30_5),
.I4(p_s1_o30_6),
.I5(p_s1_o31_0));

wire p_s2_o31_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o30_t176_z1_v0 (
.O6(p_s2_o31_2),
.O5(),
.I0(p_s1_o30_2),
.I1(p_s1_o30_3),
.I2(p_s1_o30_4),
.I3(p_s1_o30_5),
.I4(p_s1_o30_6),
.I5(p_s1_o31_0));

wire p_s2_o32_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o30_t176_z2_v0 (
.O6(p_s2_o32_0),
.O5(),
.I0(p_s1_o30_2),
.I1(p_s1_o30_3),
.I2(p_s1_o30_4),
.I3(p_s1_o30_5),
.I4(p_s1_o30_6),
.I5(p_s1_o31_0));

wire p_s2_o30_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o30_t176_z0_v1 (
.O6(p_s2_o30_5),
.O5(),
.I0(p_s1_o30_7),
.I1(p_s1_o30_8),
.I2(p_s1_o30_9),
.I3(p_s1_o30_10),
.I4(p_s1_o30_11),
.I5(p_s1_o31_1));

wire p_s2_o31_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o30_t176_z1_v1 (
.O6(p_s2_o31_3),
.O5(),
.I0(p_s1_o30_7),
.I1(p_s1_o30_8),
.I2(p_s1_o30_9),
.I3(p_s1_o30_10),
.I4(p_s1_o30_11),
.I5(p_s1_o31_1));

wire p_s2_o32_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o30_t176_z2_v1 (
.O6(p_s2_o32_1),
.O5(),
.I0(p_s1_o30_7),
.I1(p_s1_o30_8),
.I2(p_s1_o30_9),
.I3(p_s1_o30_10),
.I4(p_s1_o30_11),
.I5(p_s1_o31_1));

/////////STEP2----ORDER31////////////

wire p_s2_o31_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o31_t177_z0_v0 (
.O6(p_s2_o31_4),
.O5(),
.I0(p_s1_o31_2),
.I1(p_s1_o31_3),
.I2(p_s1_o31_4),
.I3(p_s1_o31_5),
.I4(p_s1_o31_6),
.I5(p_s1_o32_0));

wire p_s2_o32_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o31_t177_z1_v0 (
.O6(p_s2_o32_2),
.O5(),
.I0(p_s1_o31_2),
.I1(p_s1_o31_3),
.I2(p_s1_o31_4),
.I3(p_s1_o31_5),
.I4(p_s1_o31_6),
.I5(p_s1_o32_0));

wire p_s2_o33_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o31_t177_z2_v0 (
.O6(p_s2_o33_0),
.O5(),
.I0(p_s1_o31_2),
.I1(p_s1_o31_3),
.I2(p_s1_o31_4),
.I3(p_s1_o31_5),
.I4(p_s1_o31_6),
.I5(p_s1_o32_0));

wire p_s2_o31_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o31_t177_z0_v1 (
.O6(p_s2_o31_5),
.O5(),
.I0(p_s1_o31_7),
.I1(p_s1_o31_8),
.I2(p_s1_o31_9),
.I3(p_s1_o31_10),
.I4(p_s1_o31_11),
.I5(p_s1_o32_1));

wire p_s2_o32_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o31_t177_z1_v1 (
.O6(p_s2_o32_3),
.O5(),
.I0(p_s1_o31_7),
.I1(p_s1_o31_8),
.I2(p_s1_o31_9),
.I3(p_s1_o31_10),
.I4(p_s1_o31_11),
.I5(p_s1_o32_1));

wire p_s2_o33_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o31_t177_z2_v1 (
.O6(p_s2_o33_1),
.O5(),
.I0(p_s1_o31_7),
.I1(p_s1_o31_8),
.I2(p_s1_o31_9),
.I3(p_s1_o31_10),
.I4(p_s1_o31_11),
.I5(p_s1_o32_1));

/////////STEP2----ORDER32////////////

wire p_s2_o32_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o32_t178_z0_v0 (
.O6(p_s2_o32_4),
.O5(),
.I0(p_s1_o32_2),
.I1(p_s1_o32_3),
.I2(p_s1_o32_4),
.I3(p_s1_o32_5),
.I4(p_s1_o32_6),
.I5(p_s1_o33_0));

wire p_s2_o33_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o32_t178_z1_v0 (
.O6(p_s2_o33_2),
.O5(),
.I0(p_s1_o32_2),
.I1(p_s1_o32_3),
.I2(p_s1_o32_4),
.I3(p_s1_o32_5),
.I4(p_s1_o32_6),
.I5(p_s1_o33_0));

wire p_s2_o34_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o32_t178_z2_v0 (
.O6(p_s2_o34_0),
.O5(),
.I0(p_s1_o32_2),
.I1(p_s1_o32_3),
.I2(p_s1_o32_4),
.I3(p_s1_o32_5),
.I4(p_s1_o32_6),
.I5(p_s1_o33_0));

wire p_s2_o32_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o32_t178_z0_v1 (
.O6(p_s2_o32_5),
.O5(),
.I0(p_s1_o32_7),
.I1(p_s1_o32_8),
.I2(p_s1_o32_9),
.I3(p_s0_o32_15),
.I4(p_s0_o32_16),
.I5(p_s1_o33_1));

wire p_s2_o33_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o32_t178_z1_v1 (
.O6(p_s2_o33_3),
.O5(),
.I0(p_s1_o32_7),
.I1(p_s1_o32_8),
.I2(p_s1_o32_9),
.I3(p_s0_o32_15),
.I4(p_s0_o32_16),
.I5(p_s1_o33_1));

wire p_s2_o34_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o32_t178_z2_v1 (
.O6(p_s2_o34_1),
.O5(),
.I0(p_s1_o32_7),
.I1(p_s1_o32_8),
.I2(p_s1_o32_9),
.I3(p_s0_o32_15),
.I4(p_s0_o32_16),
.I5(p_s1_o33_1));

/////////STEP2----ORDER33////////////

wire p_s2_o33_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o33_t179_z0_v0 (
.O6(p_s2_o33_4),
.O5(),
.I0(p_s1_o33_2),
.I1(p_s1_o33_3),
.I2(p_s1_o33_4),
.I3(p_s1_o33_5),
.I4(p_s1_o33_6),
.I5(p_s1_o34_0));

wire p_s2_o34_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o33_t179_z1_v0 (
.O6(p_s2_o34_2),
.O5(),
.I0(p_s1_o33_2),
.I1(p_s1_o33_3),
.I2(p_s1_o33_4),
.I3(p_s1_o33_5),
.I4(p_s1_o33_6),
.I5(p_s1_o34_0));

wire p_s2_o35_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o33_t179_z2_v0 (
.O6(p_s2_o35_0),
.O5(),
.I0(p_s1_o33_2),
.I1(p_s1_o33_3),
.I2(p_s1_o33_4),
.I3(p_s1_o33_5),
.I4(p_s1_o33_6),
.I5(p_s1_o34_0));

wire p_s2_o33_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o33_t179_z0_v1 (
.O6(p_s2_o33_5),
.O5(),
.I0(p_s1_o33_7),
.I1(p_s1_o33_8),
.I2(p_s1_o33_9),
.I3(p_s1_o33_10),
.I4(p_s1_o33_11),
.I5(p_s1_o34_1));

wire p_s2_o34_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o33_t179_z1_v1 (
.O6(p_s2_o34_3),
.O5(),
.I0(p_s1_o33_7),
.I1(p_s1_o33_8),
.I2(p_s1_o33_9),
.I3(p_s1_o33_10),
.I4(p_s1_o33_11),
.I5(p_s1_o34_1));

wire p_s2_o35_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o33_t179_z2_v1 (
.O6(p_s2_o35_1),
.O5(),
.I0(p_s1_o33_7),
.I1(p_s1_o33_8),
.I2(p_s1_o33_9),
.I3(p_s1_o33_10),
.I4(p_s1_o33_11),
.I5(p_s1_o34_1));

/////////STEP2----ORDER34////////////

wire p_s2_o34_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o34_t180_z0_v0 (
.O6(p_s2_o34_4),
.O5(),
.I0(p_s1_o34_2),
.I1(p_s1_o34_3),
.I2(p_s1_o34_4),
.I3(p_s1_o34_5),
.I4(p_s1_o34_6),
.I5(p_s1_o35_0));

wire p_s2_o35_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o34_t180_z1_v0 (
.O6(p_s2_o35_2),
.O5(),
.I0(p_s1_o34_2),
.I1(p_s1_o34_3),
.I2(p_s1_o34_4),
.I3(p_s1_o34_5),
.I4(p_s1_o34_6),
.I5(p_s1_o35_0));

wire p_s2_o36_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o34_t180_z2_v0 (
.O6(p_s2_o36_0),
.O5(),
.I0(p_s1_o34_2),
.I1(p_s1_o34_3),
.I2(p_s1_o34_4),
.I3(p_s1_o34_5),
.I4(p_s1_o34_6),
.I5(p_s1_o35_0));

wire p_s2_o34_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o34_t180_z0_v1 (
.O6(p_s2_o34_5),
.O5(),
.I0(p_s1_o34_7),
.I1(p_s1_o34_8),
.I2(p_s1_o34_9),
.I3(p_s1_o34_10),
.I4(p_s1_o34_11),
.I5(p_s1_o35_1));

wire p_s2_o35_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o34_t180_z1_v1 (
.O6(p_s2_o35_3),
.O5(),
.I0(p_s1_o34_7),
.I1(p_s1_o34_8),
.I2(p_s1_o34_9),
.I3(p_s1_o34_10),
.I4(p_s1_o34_11),
.I5(p_s1_o35_1));

wire p_s2_o36_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o34_t180_z2_v1 (
.O6(p_s2_o36_1),
.O5(),
.I0(p_s1_o34_7),
.I1(p_s1_o34_8),
.I2(p_s1_o34_9),
.I3(p_s1_o34_10),
.I4(p_s1_o34_11),
.I5(p_s1_o35_1));

/////////STEP2----ORDER35////////////

wire p_s2_o35_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o35_t181_z0_v0 (
.O6(p_s2_o35_4),
.O5(),
.I0(p_s1_o35_2),
.I1(p_s1_o35_3),
.I2(p_s1_o35_4),
.I3(p_s1_o35_5),
.I4(p_s1_o35_6),
.I5(p_s1_o36_0));

wire p_s2_o36_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o35_t181_z1_v0 (
.O6(p_s2_o36_2),
.O5(),
.I0(p_s1_o35_2),
.I1(p_s1_o35_3),
.I2(p_s1_o35_4),
.I3(p_s1_o35_5),
.I4(p_s1_o35_6),
.I5(p_s1_o36_0));

wire p_s2_o37_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o35_t181_z2_v0 (
.O6(p_s2_o37_0),
.O5(),
.I0(p_s1_o35_2),
.I1(p_s1_o35_3),
.I2(p_s1_o35_4),
.I3(p_s1_o35_5),
.I4(p_s1_o35_6),
.I5(p_s1_o36_0));

wire p_s2_o35_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o35_t181_z0_v1 (
.O6(p_s2_o35_5),
.O5(),
.I0(p_s1_o35_7),
.I1(p_s1_o35_8),
.I2(p_s1_o35_9),
.I3(p_s1_o35_10),
.I4(p_s1_o35_11),
.I5(p_s1_o36_1));

wire p_s2_o36_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o35_t181_z1_v1 (
.O6(p_s2_o36_3),
.O5(),
.I0(p_s1_o35_7),
.I1(p_s1_o35_8),
.I2(p_s1_o35_9),
.I3(p_s1_o35_10),
.I4(p_s1_o35_11),
.I5(p_s1_o36_1));

wire p_s2_o37_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o35_t181_z2_v1 (
.O6(p_s2_o37_1),
.O5(),
.I0(p_s1_o35_7),
.I1(p_s1_o35_8),
.I2(p_s1_o35_9),
.I3(p_s1_o35_10),
.I4(p_s1_o35_11),
.I5(p_s1_o36_1));

/////////STEP2----ORDER36////////////

wire p_s2_o36_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o36_t182_z0_v0 (
.O6(p_s2_o36_4),
.O5(),
.I0(p_s1_o36_2),
.I1(p_s1_o36_3),
.I2(p_s1_o36_4),
.I3(p_s1_o36_5),
.I4(p_s1_o36_6),
.I5(p_s1_o37_0));

wire p_s2_o37_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o36_t182_z1_v0 (
.O6(p_s2_o37_2),
.O5(),
.I0(p_s1_o36_2),
.I1(p_s1_o36_3),
.I2(p_s1_o36_4),
.I3(p_s1_o36_5),
.I4(p_s1_o36_6),
.I5(p_s1_o37_0));

wire p_s2_o38_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o36_t182_z2_v0 (
.O6(p_s2_o38_0),
.O5(),
.I0(p_s1_o36_2),
.I1(p_s1_o36_3),
.I2(p_s1_o36_4),
.I3(p_s1_o36_5),
.I4(p_s1_o36_6),
.I5(p_s1_o37_0));

wire p_s2_o36_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o36_t182_z0_v1 (
.O6(p_s2_o36_5),
.O5(),
.I0(p_s1_o36_7),
.I1(p_s1_o36_8),
.I2(p_s1_o36_9),
.I3(p_s1_o36_10),
.I4(p_s1_o36_11),
.I5(p_s1_o37_1));

wire p_s2_o37_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o36_t182_z1_v1 (
.O6(p_s2_o37_3),
.O5(),
.I0(p_s1_o36_7),
.I1(p_s1_o36_8),
.I2(p_s1_o36_9),
.I3(p_s1_o36_10),
.I4(p_s1_o36_11),
.I5(p_s1_o37_1));

wire p_s2_o38_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o36_t182_z2_v1 (
.O6(p_s2_o38_1),
.O5(),
.I0(p_s1_o36_7),
.I1(p_s1_o36_8),
.I2(p_s1_o36_9),
.I3(p_s1_o36_10),
.I4(p_s1_o36_11),
.I5(p_s1_o37_1));

/////////STEP2----ORDER37////////////

wire p_s2_o37_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o37_t183_z0_v0 (
.O6(p_s2_o37_4),
.O5(),
.I0(p_s1_o37_2),
.I1(p_s1_o37_3),
.I2(p_s1_o37_4),
.I3(p_s1_o37_5),
.I4(p_s1_o37_6),
.I5(p_s1_o38_0));

wire p_s2_o38_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o37_t183_z1_v0 (
.O6(p_s2_o38_2),
.O5(),
.I0(p_s1_o37_2),
.I1(p_s1_o37_3),
.I2(p_s1_o37_4),
.I3(p_s1_o37_5),
.I4(p_s1_o37_6),
.I5(p_s1_o38_0));

wire p_s2_o39_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o37_t183_z2_v0 (
.O6(p_s2_o39_0),
.O5(),
.I0(p_s1_o37_2),
.I1(p_s1_o37_3),
.I2(p_s1_o37_4),
.I3(p_s1_o37_5),
.I4(p_s1_o37_6),
.I5(p_s1_o38_0));

wire p_s2_o37_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o37_t183_z0_v1 (
.O6(p_s2_o37_5),
.O5(),
.I0(p_s1_o37_7),
.I1(p_s1_o37_8),
.I2(p_s1_o37_9),
.I3(p_s1_o37_10),
.I4(p_s1_o37_11),
.I5(p_s1_o38_1));

wire p_s2_o38_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o37_t183_z1_v1 (
.O6(p_s2_o38_3),
.O5(),
.I0(p_s1_o37_7),
.I1(p_s1_o37_8),
.I2(p_s1_o37_9),
.I3(p_s1_o37_10),
.I4(p_s1_o37_11),
.I5(p_s1_o38_1));

wire p_s2_o39_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o37_t183_z2_v1 (
.O6(p_s2_o39_1),
.O5(),
.I0(p_s1_o37_7),
.I1(p_s1_o37_8),
.I2(p_s1_o37_9),
.I3(p_s1_o37_10),
.I4(p_s1_o37_11),
.I5(p_s1_o38_1));

/////////STEP2----ORDER38////////////

wire p_s2_o38_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o38_t184_z0_v0 (
.O6(p_s2_o38_4),
.O5(),
.I0(p_s1_o38_2),
.I1(p_s1_o38_3),
.I2(p_s1_o38_4),
.I3(p_s1_o38_5),
.I4(p_s1_o38_6),
.I5(p_s1_o39_0));

wire p_s2_o39_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o38_t184_z1_v0 (
.O6(p_s2_o39_2),
.O5(),
.I0(p_s1_o38_2),
.I1(p_s1_o38_3),
.I2(p_s1_o38_4),
.I3(p_s1_o38_5),
.I4(p_s1_o38_6),
.I5(p_s1_o39_0));

wire p_s2_o40_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o38_t184_z2_v0 (
.O6(p_s2_o40_0),
.O5(),
.I0(p_s1_o38_2),
.I1(p_s1_o38_3),
.I2(p_s1_o38_4),
.I3(p_s1_o38_5),
.I4(p_s1_o38_6),
.I5(p_s1_o39_0));

wire p_s2_o38_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o38_t184_z0_v1 (
.O6(p_s2_o38_5),
.O5(),
.I0(p_s1_o38_7),
.I1(p_s1_o38_8),
.I2(p_s1_o38_9),
.I3(p_s1_o38_10),
.I4(p_s1_o38_11),
.I5(p_s1_o39_1));

wire p_s2_o39_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o38_t184_z1_v1 (
.O6(p_s2_o39_3),
.O5(),
.I0(p_s1_o38_7),
.I1(p_s1_o38_8),
.I2(p_s1_o38_9),
.I3(p_s1_o38_10),
.I4(p_s1_o38_11),
.I5(p_s1_o39_1));

wire p_s2_o40_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o38_t184_z2_v1 (
.O6(p_s2_o40_1),
.O5(),
.I0(p_s1_o38_7),
.I1(p_s1_o38_8),
.I2(p_s1_o38_9),
.I3(p_s1_o38_10),
.I4(p_s1_o38_11),
.I5(p_s1_o39_1));

/////////STEP2----ORDER39////////////

wire p_s2_o39_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o39_t185_z0_v0 (
.O6(p_s2_o39_4),
.O5(),
.I0(p_s1_o39_2),
.I1(p_s1_o39_3),
.I2(p_s1_o39_4),
.I3(p_s1_o39_5),
.I4(p_s1_o39_6),
.I5(p_s1_o40_0));

wire p_s2_o40_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o39_t185_z1_v0 (
.O6(p_s2_o40_2),
.O5(),
.I0(p_s1_o39_2),
.I1(p_s1_o39_3),
.I2(p_s1_o39_4),
.I3(p_s1_o39_5),
.I4(p_s1_o39_6),
.I5(p_s1_o40_0));

wire p_s2_o41_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o39_t185_z2_v0 (
.O6(p_s2_o41_0),
.O5(),
.I0(p_s1_o39_2),
.I1(p_s1_o39_3),
.I2(p_s1_o39_4),
.I3(p_s1_o39_5),
.I4(p_s1_o39_6),
.I5(p_s1_o40_0));

wire p_s2_o39_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o39_t185_z0_v1 (
.O6(p_s2_o39_5),
.O5(),
.I0(p_s1_o39_7),
.I1(p_s1_o39_8),
.I2(p_s1_o39_9),
.I3(p_s1_o39_10),
.I4(p_s1_o39_11),
.I5(p_s1_o40_1));

wire p_s2_o40_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o39_t185_z1_v1 (
.O6(p_s2_o40_3),
.O5(),
.I0(p_s1_o39_7),
.I1(p_s1_o39_8),
.I2(p_s1_o39_9),
.I3(p_s1_o39_10),
.I4(p_s1_o39_11),
.I5(p_s1_o40_1));

wire p_s2_o41_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o39_t185_z2_v1 (
.O6(p_s2_o41_1),
.O5(),
.I0(p_s1_o39_7),
.I1(p_s1_o39_8),
.I2(p_s1_o39_9),
.I3(p_s1_o39_10),
.I4(p_s1_o39_11),
.I5(p_s1_o40_1));

/////////STEP2----ORDER40////////////

wire p_s2_o40_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o40_t186_z0_v0 (
.O6(p_s2_o40_4),
.O5(),
.I0(p_s1_o40_2),
.I1(p_s1_o40_3),
.I2(p_s1_o40_4),
.I3(p_s1_o40_5),
.I4(p_s1_o40_6),
.I5(p_s1_o41_0));

wire p_s2_o41_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o40_t186_z1_v0 (
.O6(p_s2_o41_2),
.O5(),
.I0(p_s1_o40_2),
.I1(p_s1_o40_3),
.I2(p_s1_o40_4),
.I3(p_s1_o40_5),
.I4(p_s1_o40_6),
.I5(p_s1_o41_0));

wire p_s2_o42_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o40_t186_z2_v0 (
.O6(p_s2_o42_0),
.O5(),
.I0(p_s1_o40_2),
.I1(p_s1_o40_3),
.I2(p_s1_o40_4),
.I3(p_s1_o40_5),
.I4(p_s1_o40_6),
.I5(p_s1_o41_0));

wire p_s2_o40_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o40_t186_z0_v1 (
.O6(p_s2_o40_5),
.O5(),
.I0(p_s1_o40_7),
.I1(p_s1_o40_8),
.I2(p_s1_o40_9),
.I3(p_s1_o40_10),
.I4(p_s1_o40_11),
.I5(p_s1_o41_1));

wire p_s2_o41_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o40_t186_z1_v1 (
.O6(p_s2_o41_3),
.O5(),
.I0(p_s1_o40_7),
.I1(p_s1_o40_8),
.I2(p_s1_o40_9),
.I3(p_s1_o40_10),
.I4(p_s1_o40_11),
.I5(p_s1_o41_1));

wire p_s2_o42_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o40_t186_z2_v1 (
.O6(p_s2_o42_1),
.O5(),
.I0(p_s1_o40_7),
.I1(p_s1_o40_8),
.I2(p_s1_o40_9),
.I3(p_s1_o40_10),
.I4(p_s1_o40_11),
.I5(p_s1_o41_1));

/////////STEP2----ORDER41////////////

wire p_s2_o41_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o41_t187_z0_v0 (
.O6(p_s2_o41_4),
.O5(),
.I0(p_s1_o41_2),
.I1(p_s1_o41_3),
.I2(p_s1_o41_4),
.I3(p_s1_o41_5),
.I4(p_s1_o41_6),
.I5(p_s1_o42_0));

wire p_s2_o42_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o41_t187_z1_v0 (
.O6(p_s2_o42_2),
.O5(),
.I0(p_s1_o41_2),
.I1(p_s1_o41_3),
.I2(p_s1_o41_4),
.I3(p_s1_o41_5),
.I4(p_s1_o41_6),
.I5(p_s1_o42_0));

wire p_s2_o43_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o41_t187_z2_v0 (
.O6(p_s2_o43_0),
.O5(),
.I0(p_s1_o41_2),
.I1(p_s1_o41_3),
.I2(p_s1_o41_4),
.I3(p_s1_o41_5),
.I4(p_s1_o41_6),
.I5(p_s1_o42_0));

wire p_s2_o41_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o41_t187_z0_v1 (
.O6(p_s2_o41_5),
.O5(),
.I0(p_s1_o41_7),
.I1(p_s1_o41_8),
.I2(p_s1_o41_9),
.I3(p_s1_o41_10),
.I4(p_s1_o41_11),
.I5(p_s1_o42_1));

wire p_s2_o42_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o41_t187_z1_v1 (
.O6(p_s2_o42_3),
.O5(),
.I0(p_s1_o41_7),
.I1(p_s1_o41_8),
.I2(p_s1_o41_9),
.I3(p_s1_o41_10),
.I4(p_s1_o41_11),
.I5(p_s1_o42_1));

wire p_s2_o43_1;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o41_t187_z2_v1 (
.O6(p_s2_o43_1),
.O5(),
.I0(p_s1_o41_7),
.I1(p_s1_o41_8),
.I2(p_s1_o41_9),
.I3(p_s1_o41_10),
.I4(p_s1_o41_11),
.I5(p_s1_o42_1));

/////////STEP2----ORDER42////////////

wire p_s2_o42_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o42_t188_z0_v0 (
.O6(p_s2_o42_4),
.O5(),
.I0(p_s1_o42_2),
.I1(p_s1_o42_3),
.I2(p_s1_o42_4),
.I3(p_s1_o42_5),
.I4(p_s1_o42_6),
.I5(p_s1_o43_0));

wire p_s2_o43_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o42_t188_z1_v0 (
.O6(p_s2_o43_2),
.O5(),
.I0(p_s1_o42_2),
.I1(p_s1_o42_3),
.I2(p_s1_o42_4),
.I3(p_s1_o42_5),
.I4(p_s1_o42_6),
.I5(p_s1_o43_0));

wire p_s2_o44_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o42_t188_z2_v0 (
.O6(p_s2_o44_0),
.O5(),
.I0(p_s1_o42_2),
.I1(p_s1_o42_3),
.I2(p_s1_o42_4),
.I3(p_s1_o42_5),
.I4(p_s1_o42_6),
.I5(p_s1_o43_0));

wire p_s2_o43_3;
wire p_s2_o42_5;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s2_o42_t193_z0_v0 (
.O6(p_s2_o43_3),
.O5(p_s2_o42_5),
.I0(p_s1_o42_7),
.I1(p_s1_o42_8),
.I2(p_s1_o42_9),
.I3(p_s1_o43_1),
.I4(p_s1_o43_2),
.I5(1'b1));

wire p_s2_o44_1;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s2_o42_t193_z1_v0 (
.O6(p_s2_o44_1),
.O5(),
.I0(p_s1_o42_7),
.I1(p_s1_o42_8),
.I2(p_s1_o42_9),
.I3(p_s1_o43_1),
.I4(p_s1_o43_2),
.I5(1'b1));

/////////STEP2----ORDER43////////////

wire p_s2_o44_2;
wire p_s2_o43_4;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o43_t133_z0_v0 (
.O6(p_s2_o44_2),
.O5(p_s2_o43_4),
.I0(a[15]),
.I1(b[31]),
.I2(p_s1_o43_3),
.I3(p_s1_o43_4),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o43_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o43_t189_z0_v0 (
.O6(p_s2_o43_5),
.O5(),
.I0(p_s1_o43_5),
.I1(p_s1_o43_6),
.I2(p_s1_o43_7),
.I3(p_s1_o43_8),
.I4(p_s1_o43_9),
.I5(p_s1_o44_0));

wire p_s2_o44_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o43_t189_z1_v0 (
.O6(p_s2_o44_3),
.O5(),
.I0(p_s1_o43_5),
.I1(p_s1_o43_6),
.I2(p_s1_o43_7),
.I3(p_s1_o43_8),
.I4(p_s1_o43_9),
.I5(p_s1_o44_0));

wire p_s2_o45_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o43_t189_z2_v0 (
.O6(p_s2_o45_0),
.O5(),
.I0(p_s1_o43_5),
.I1(p_s1_o43_6),
.I2(p_s1_o43_7),
.I3(p_s1_o43_8),
.I4(p_s1_o43_9),
.I5(p_s1_o44_0));

/////////STEP2----ORDER44////////////

wire p_s2_o45_1;
wire p_s2_o44_4;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s2_o44_t128_z0_v0 (
.O6(p_s2_o45_1),
.O5(p_s2_o44_4),
.I0(p_s1_o44_1),
.I1(p_s1_o44_2),
.I2(p_s1_o44_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o44_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o44_t190_z0_v0 (
.O6(p_s2_o44_5),
.O5(),
.I0(p_s1_o44_4),
.I1(p_s1_o44_5),
.I2(p_s1_o44_6),
.I3(p_s1_o44_7),
.I4(p_s1_o44_8),
.I5(p_s1_o45_0));

wire p_s2_o45_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o44_t190_z1_v0 (
.O6(p_s2_o45_2),
.O5(),
.I0(p_s1_o44_4),
.I1(p_s1_o44_5),
.I2(p_s1_o44_6),
.I3(p_s1_o44_7),
.I4(p_s1_o44_8),
.I5(p_s1_o45_0));

wire p_s2_o46_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o44_t190_z2_v0 (
.O6(p_s2_o46_0),
.O5(),
.I0(p_s1_o44_4),
.I1(p_s1_o44_5),
.I2(p_s1_o44_6),
.I3(p_s1_o44_7),
.I4(p_s1_o44_8),
.I5(p_s1_o45_0));

/////////STEP2----ORDER45////////////

wire p_s2_o46_1;
wire p_s2_o45_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o45_t145_z0_v0 (
.O6(p_s2_o46_1),
.O5(p_s2_o45_3),
.I0(a[20]),
.I1(b[28]),
.I2(a[19]),
.I3(b[29]),
.I4(p_s1_o45_1),
.I5(1'b1));

wire p_s2_o46_2;
wire p_s2_o45_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o45_t145_z0_v1 (
.O6(p_s2_o46_2),
.O5(p_s2_o45_4),
.I0(a[18]),
.I1(b[30]),
.I2(a[17]),
.I3(b[31]),
.I4(p_s1_o45_2),
.I5(1'b1));

wire p_s2_o45_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o45_t191_z0_v0 (
.O6(p_s2_o45_5),
.O5(),
.I0(p_s1_o45_3),
.I1(p_s1_o45_4),
.I2(p_s1_o45_5),
.I3(p_s1_o45_6),
.I4(p_s1_o45_7),
.I5(p_s1_o46_0));

wire p_s2_o46_3;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o45_t191_z1_v0 (
.O6(p_s2_o46_3),
.O5(),
.I0(p_s1_o45_3),
.I1(p_s1_o45_4),
.I2(p_s1_o45_5),
.I3(p_s1_o45_6),
.I4(p_s1_o45_7),
.I5(p_s1_o46_0));

wire p_s2_o47_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o45_t191_z2_v0 (
.O6(p_s2_o47_0),
.O5(),
.I0(p_s1_o45_3),
.I1(p_s1_o45_4),
.I2(p_s1_o45_5),
.I3(p_s1_o45_6),
.I4(p_s1_o45_7),
.I5(p_s1_o46_0));

/////////STEP2----ORDER46////////////

wire p_s2_o47_1;
wire p_s2_o46_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o46_t146_z0_v0 (
.O6(p_s2_o47_1),
.O5(p_s2_o46_4),
.I0(a[19]),
.I1(b[30]),
.I2(a[18]),
.I3(b[31]),
.I4(p_s1_o46_1),
.I5(1'b1));

wire p_s2_o46_5;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o46_t192_z0_v0 (
.O6(p_s2_o46_5),
.O5(),
.I0(p_s1_o46_2),
.I1(p_s1_o46_3),
.I2(p_s1_o46_4),
.I3(p_s1_o46_5),
.I4(p_s1_o46_6),
.I5(p_s1_o47_0));

wire p_s2_o47_2;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o46_t192_z1_v0 (
.O6(p_s2_o47_2),
.O5(),
.I0(p_s1_o46_2),
.I1(p_s1_o46_3),
.I2(p_s1_o46_4),
.I3(p_s1_o46_5),
.I4(p_s1_o46_6),
.I5(p_s1_o47_0));

wire p_s2_o48_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o46_t192_z2_v0 (
.O6(p_s2_o48_0),
.O5(),
.I0(p_s1_o46_2),
.I1(p_s1_o46_3),
.I2(p_s1_o46_4),
.I3(p_s1_o46_5),
.I4(p_s1_o46_6),
.I5(p_s1_o47_0));

/////////STEP2----ORDER47////////////

wire p_s2_o48_1;
wire p_s2_o47_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o47_t147_z0_v0 (
.O6(p_s2_o48_1),
.O5(p_s2_o47_3),
.I0(a[22]),
.I1(b[28]),
.I2(a[21]),
.I3(b[29]),
.I4(p_s1_o47_1),
.I5(1'b1));

wire p_s2_o48_2;
wire p_s2_o47_4;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s2_o47_t194_z0_v0 (
.O6(p_s2_o48_2),
.O5(p_s2_o47_4),
.I0(p_s1_o47_2),
.I1(p_s1_o47_3),
.I2(p_s1_o47_4),
.I3(p_s1_o48_0),
.I4(p_s1_o48_1),
.I5(1'b1));

wire p_s2_o49_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s2_o47_t194_z1_v0 (
.O6(p_s2_o49_0),
.O5(),
.I0(p_s1_o47_2),
.I1(p_s1_o47_3),
.I2(p_s1_o47_4),
.I3(p_s1_o48_0),
.I4(p_s1_o48_1),
.I5(1'b1));

/////////STEP2----ORDER48////////////

wire p_s2_o49_1;
wire p_s2_o48_3;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s2_o48_t129_z0_v0 (
.O6(p_s2_o49_1),
.O5(p_s2_o48_3),
.I0(p_s1_o48_2),
.I1(p_s1_o48_3),
.I2(p_s1_o48_4),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP2----ORDER49////////////

wire p_s2_o50_0;
wire p_s2_o49_2;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o49_t134_z0_v0 (
.O6(p_s2_o50_0),
.O5(p_s2_o49_2),
.I0(a[27]),
.I1(b[25]),
.I2(p_s1_o49_0),
.I3(p_s1_o49_1),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o50_1;
wire p_s2_o49_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o49_t148_z0_v0 (
.O6(p_s2_o50_1),
.O5(p_s2_o49_3),
.I0(a[26]),
.I1(b[26]),
.I2(a[25]),
.I3(b[27]),
.I4(p_s1_o49_2),
.I5(1'b1));

wire p_s2_o50_2;
wire p_s2_o49_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o49_t148_z0_v1 (
.O6(p_s2_o50_2),
.O5(p_s2_o49_4),
.I0(a[24]),
.I1(b[28]),
.I2(a[23]),
.I3(b[29]),
.I4(p_s1_o49_3),
.I5(1'b1));

wire p_s2_o50_3;
wire p_s2_o49_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o49_t148_z0_v2 (
.O6(p_s2_o50_3),
.O5(p_s2_o49_5),
.I0(a[22]),
.I1(b[30]),
.I2(a[21]),
.I3(b[31]),
.I4(p_s1_o49_4),
.I5(1'b1));

/////////STEP2----ORDER50////////////

wire p_s2_o51_0;
wire p_s2_o50_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o50_t149_z0_v0 (
.O6(p_s2_o51_0),
.O5(p_s2_o50_4),
.I0(a[28]),
.I1(b[25]),
.I2(a[27]),
.I3(b[26]),
.I4(p_s1_o50_0),
.I5(1'b1));

wire p_s2_o51_1;
wire p_s2_o50_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o50_t149_z0_v1 (
.O6(p_s2_o51_1),
.O5(p_s2_o50_5),
.I0(a[26]),
.I1(b[27]),
.I2(a[25]),
.I3(b[28]),
.I4(p_s1_o50_1),
.I5(1'b1));

wire p_s2_o51_2;
wire p_s2_o50_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o50_t149_z0_v2 (
.O6(p_s2_o51_2),
.O5(p_s2_o50_6),
.I0(a[24]),
.I1(b[29]),
.I2(a[23]),
.I3(b[30]),
.I4(p_s0_o50_0),
.I5(1'b1));

/////////STEP2----ORDER51////////////

wire p_s2_o52_0;
wire p_s2_o51_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o51_t150_z0_v0 (
.O6(p_s2_o52_0),
.O5(p_s2_o51_3),
.I0(a[24]),
.I1(b[30]),
.I2(a[23]),
.I3(b[31]),
.I4(p_s1_o51_0),
.I5(1'b1));

/////////STEP2----ORDER52////////////

wire p_s2_o53_0;
wire p_s2_o52_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o52_t151_z0_v0 (
.O6(p_s2_o53_0),
.O5(p_s2_o52_1),
.I0(a[29]),
.I1(b[26]),
.I2(a[28]),
.I3(b[27]),
.I4(p_s1_o52_0),
.I5(1'b1));

wire p_s2_o53_1;
wire p_s2_o52_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o52_t151_z0_v1 (
.O6(p_s2_o53_1),
.O5(p_s2_o52_2),
.I0(a[27]),
.I1(b[28]),
.I2(a[26]),
.I3(b[29]),
.I4(p_s1_o52_1),
.I5(1'b1));

wire p_s2_o53_2;
wire p_s2_o52_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o52_t151_z0_v2 (
.O6(p_s2_o53_2),
.O5(p_s2_o52_3),
.I0(a[25]),
.I1(b[30]),
.I2(a[24]),
.I3(b[31]),
.I4(p_s1_o52_2),
.I5(1'b1));

/////////STEP2----ORDER53////////////

wire p_s2_o54_0;
wire p_s2_o53_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o53_t152_z0_v0 (
.O6(p_s2_o54_0),
.O5(p_s2_o53_3),
.I0(a[31]),
.I1(b[25]),
.I2(a[30]),
.I3(b[26]),
.I4(p_s1_o53_0),
.I5(1'b1));

/////////STEP2----ORDER54////////////

/////////STEP2----ORDER55////////////

wire p_s2_o56_0;
wire p_s2_o55_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o55_t153_z0_v0 (
.O6(p_s2_o56_0),
.O5(p_s2_o55_0),
.I0(a[29]),
.I1(b[29]),
.I2(a[28]),
.I3(b[30]),
.I4(p_s1_o55_0),
.I5(1'b1));

/////////STEP2----ORDER56////////////

wire p_s2_o57_0;
wire p_s2_o56_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o56_t154_z0_v0 (
.O6(p_s2_o57_0),
.O5(p_s2_o56_1),
.I0(a[31]),
.I1(b[28]),
.I2(a[30]),
.I3(b[29]),
.I4(p_s1_o56_0),
.I5(1'b1));

/////////STEP2----ORDER57////////////

/////////STEP2----ORDER58////////////

/////////STEP2----ORDER59////////////

/////////STEP3----ORDER0////////////

/////////STEP3----ORDER1////////////

/////////STEP3----ORDER2////////////

wire p_s3_o3_0;
wire p_s3_o2_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o2_t213_z0_v0 (
.O6(p_s3_o3_0),
.O5(p_s3_o2_0),
.I0(a[3]),
.I1(b[2]),
.I2(a[2]),
.I3(b[3]),
.I4(p_s2_o2_0),
.I5(1'b1));

wire p_s3_o3_1;
wire p_s3_o2_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o2_t213_z0_v1 (
.O6(p_s3_o3_1),
.O5(p_s3_o2_1),
.I0(a[1]),
.I1(b[4]),
.I2(a[0]),
.I3(b[5]),
.I4(p_s2_o2_1),
.I5(1'b1));

/////////STEP3----ORDER3////////////

/////////STEP3----ORDER4////////////

wire p_s3_o5_0;
wire p_s3_o4_0;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o4_t206_z0_v0 (
.O6(p_s3_o5_0),
.O5(p_s3_o4_0),
.I0(a[0]),
.I1(b[7]),
.I2(p_s2_o4_0),
.I3(p_s1_o4_0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER5////////////

wire p_s3_o6_0;
wire p_s3_o5_1;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o5_t207_z0_v0 (
.O6(p_s3_o6_0),
.O5(p_s3_o5_1),
.I0(a[0]),
.I1(b[8]),
.I2(p_s2_o5_0),
.I3(p_s2_o5_1),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER6////////////

wire p_s3_o7_0;
wire p_s3_o6_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o6_t214_z0_v0 (
.O6(p_s3_o7_0),
.O5(p_s3_o6_1),
.I0(a[7]),
.I1(b[2]),
.I2(a[6]),
.I3(b[3]),
.I4(p_s2_o6_0),
.I5(1'b1));

wire p_s3_o7_1;
wire p_s3_o6_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o6_t214_z0_v1 (
.O6(p_s3_o7_1),
.O5(p_s3_o6_2),
.I0(a[5]),
.I1(b[4]),
.I2(a[4]),
.I3(b[5]),
.I4(p_s2_o6_1),
.I5(1'b1));

wire p_s3_o7_2;
wire p_s3_o6_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o6_t214_z0_v2 (
.O6(p_s3_o7_2),
.O5(p_s3_o6_3),
.I0(a[3]),
.I1(b[6]),
.I2(a[2]),
.I3(b[7]),
.I4(p_s2_o6_2),
.I5(1'b1));

wire p_s3_o7_3;
wire p_s3_o6_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o6_t214_z0_v3 (
.O6(p_s3_o7_3),
.O5(p_s3_o6_4),
.I0(a[1]),
.I1(b[8]),
.I2(a[0]),
.I3(b[9]),
.I4(p_s2_o6_3),
.I5(1'b1));

/////////STEP3----ORDER7////////////

/////////STEP3----ORDER8////////////

wire p_s3_o8_0;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o8_t224_z0_v0 (
.O6(p_s3_o8_0),
.O5(),
.I0(p_s2_o8_0),
.I1(p_s2_o8_1),
.I2(p_s2_o8_2),
.I3(p_s2_o8_3),
.I4(p_s2_o8_4),
.I5(p_s2_o9_0));

wire p_s3_o9_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o8_t224_z1_v0 (
.O6(p_s3_o9_0),
.O5(),
.I0(p_s2_o8_0),
.I1(p_s2_o8_1),
.I2(p_s2_o8_2),
.I3(p_s2_o8_3),
.I4(p_s2_o8_4),
.I5(p_s2_o9_0));

wire p_s3_o10_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o8_t224_z2_v0 (
.O6(p_s3_o10_0),
.O5(),
.I0(p_s2_o8_0),
.I1(p_s2_o8_1),
.I2(p_s2_o8_2),
.I3(p_s2_o8_3),
.I4(p_s2_o8_4),
.I5(p_s2_o9_0));

/////////STEP3----ORDER9////////////

wire p_s3_o10_1;
wire p_s3_o9_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o9_t195_z0_v0 (
.O6(p_s3_o10_1),
.O5(p_s3_o9_1),
.I0(p_s2_o9_1),
.I1(p_s2_o9_2),
.I2(p_s2_o9_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o10_2;
wire p_s3_o9_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o9_t215_z0_v0 (
.O6(p_s3_o10_2),
.O5(p_s3_o9_2),
.I0(a[1]),
.I1(b[11]),
.I2(a[0]),
.I3(b[12]),
.I4(p_s2_o9_4),
.I5(1'b1));

/////////STEP3----ORDER10////////////

wire p_s3_o10_3;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o10_t225_z0_v0 (
.O6(p_s3_o10_3),
.O5(),
.I0(p_s2_o10_0),
.I1(p_s2_o10_1),
.I2(p_s2_o10_2),
.I3(p_s2_o10_3),
.I4(p_s2_o10_4),
.I5(p_s2_o11_0));

wire p_s3_o11_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o10_t225_z1_v0 (
.O6(p_s3_o11_0),
.O5(),
.I0(p_s2_o10_0),
.I1(p_s2_o10_1),
.I2(p_s2_o10_2),
.I3(p_s2_o10_3),
.I4(p_s2_o10_4),
.I5(p_s2_o11_0));

wire p_s3_o12_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o10_t225_z2_v0 (
.O6(p_s3_o12_0),
.O5(),
.I0(p_s2_o10_0),
.I1(p_s2_o10_1),
.I2(p_s2_o10_2),
.I3(p_s2_o10_3),
.I4(p_s2_o10_4),
.I5(p_s2_o11_0));

/////////STEP3----ORDER11////////////

wire p_s3_o12_1;
wire p_s3_o11_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o11_t196_z0_v0 (
.O6(p_s3_o12_1),
.O5(p_s3_o11_1),
.I0(p_s2_o11_1),
.I1(p_s2_o11_2),
.I2(p_s2_o11_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER12////////////

wire p_s3_o12_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o12_t226_z0_v0 (
.O6(p_s3_o12_2),
.O5(),
.I0(p_s2_o12_0),
.I1(p_s2_o12_1),
.I2(p_s2_o12_2),
.I3(p_s2_o12_3),
.I4(p_s2_o12_4),
.I5(p_s2_o13_0));

wire p_s3_o13_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o12_t226_z1_v0 (
.O6(p_s3_o13_0),
.O5(),
.I0(p_s2_o12_0),
.I1(p_s2_o12_1),
.I2(p_s2_o12_2),
.I3(p_s2_o12_3),
.I4(p_s2_o12_4),
.I5(p_s2_o13_0));

wire p_s3_o14_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o12_t226_z2_v0 (
.O6(p_s3_o14_0),
.O5(),
.I0(p_s2_o12_0),
.I1(p_s2_o12_1),
.I2(p_s2_o12_2),
.I3(p_s2_o12_3),
.I4(p_s2_o12_4),
.I5(p_s2_o13_0));

/////////STEP3----ORDER13////////////

wire p_s3_o13_1;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s3_o13_t219_z0_v0 (
.O6(p_s3_o13_1),
.O5(),
.I0(p_s2_o13_1),
.I1(p_s2_o13_2),
.I2(p_s2_o13_3),
.I3(p_s2_o13_4),
.I4(p_s2_o13_5),
.I5(p_s2_o13_6));

wire p_s3_o14_1;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s3_o13_t219_z1_v0 (
.O6(p_s3_o14_1),
.O5(),
.I0(p_s2_o13_1),
.I1(p_s2_o13_2),
.I2(p_s2_o13_3),
.I3(p_s2_o13_4),
.I4(p_s2_o13_5),
.I5(p_s2_o13_6));

wire p_s3_o15_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s3_o13_t219_z2_v0 (
.O6(p_s3_o15_0),
.O5(),
.I0(p_s2_o13_1),
.I1(p_s2_o13_2),
.I2(p_s2_o13_3),
.I3(p_s2_o13_4),
.I4(p_s2_o13_5),
.I5(p_s2_o13_6));

/////////STEP3----ORDER14////////////

/////////STEP3----ORDER15////////////

/////////STEP3----ORDER16////////////

wire p_s3_o16_0;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s3_o16_t220_z0_v0 (
.O6(p_s3_o16_0),
.O5(),
.I0(p_s2_o16_0),
.I1(p_s2_o16_1),
.I2(p_s2_o16_2),
.I3(p_s2_o16_3),
.I4(p_s2_o16_4),
.I5(p_s2_o16_5));

wire p_s3_o17_0;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s3_o16_t220_z1_v0 (
.O6(p_s3_o17_0),
.O5(),
.I0(p_s2_o16_0),
.I1(p_s2_o16_1),
.I2(p_s2_o16_2),
.I3(p_s2_o16_3),
.I4(p_s2_o16_4),
.I5(p_s2_o16_5));

wire p_s3_o18_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s3_o16_t220_z2_v0 (
.O6(p_s3_o18_0),
.O5(),
.I0(p_s2_o16_0),
.I1(p_s2_o16_1),
.I2(p_s2_o16_2),
.I3(p_s2_o16_3),
.I4(p_s2_o16_4),
.I5(p_s2_o16_5));

/////////STEP3----ORDER17////////////

wire p_s3_o18_1;
wire p_s3_o17_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o17_t197_z0_v0 (
.O6(p_s3_o18_1),
.O5(p_s3_o17_1),
.I0(p_s2_o17_0),
.I1(p_s2_o17_1),
.I2(p_s2_o17_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o18_2;
wire p_s3_o17_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o17_t197_z0_v1 (
.O6(p_s3_o18_2),
.O5(p_s3_o17_2),
.I0(p_s2_o17_3),
.I1(p_s2_o17_4),
.I2(p_s2_o17_5),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER18////////////

wire p_s3_o18_3;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o18_t227_z0_v0 (
.O6(p_s3_o18_3),
.O5(),
.I0(p_s2_o18_0),
.I1(p_s2_o18_1),
.I2(p_s2_o18_2),
.I3(p_s2_o18_3),
.I4(p_s2_o18_4),
.I5(p_s2_o19_0));

wire p_s3_o19_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o18_t227_z1_v0 (
.O6(p_s3_o19_0),
.O5(),
.I0(p_s2_o18_0),
.I1(p_s2_o18_1),
.I2(p_s2_o18_2),
.I3(p_s2_o18_3),
.I4(p_s2_o18_4),
.I5(p_s2_o19_0));

wire p_s3_o20_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o18_t227_z2_v0 (
.O6(p_s3_o20_0),
.O5(),
.I0(p_s2_o18_0),
.I1(p_s2_o18_1),
.I2(p_s2_o18_2),
.I3(p_s2_o18_3),
.I4(p_s2_o18_4),
.I5(p_s2_o19_0));

/////////STEP3----ORDER19////////////

wire p_s3_o19_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o19_t228_z0_v0 (
.O6(p_s3_o19_1),
.O5(),
.I0(p_s2_o19_1),
.I1(p_s2_o19_2),
.I2(p_s2_o19_3),
.I3(p_s2_o19_4),
.I4(p_s2_o19_5),
.I5(p_s2_o20_0));

wire p_s3_o20_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o19_t228_z1_v0 (
.O6(p_s3_o20_1),
.O5(),
.I0(p_s2_o19_1),
.I1(p_s2_o19_2),
.I2(p_s2_o19_3),
.I3(p_s2_o19_4),
.I4(p_s2_o19_5),
.I5(p_s2_o20_0));

wire p_s3_o21_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o19_t228_z2_v0 (
.O6(p_s3_o21_0),
.O5(),
.I0(p_s2_o19_1),
.I1(p_s2_o19_2),
.I2(p_s2_o19_3),
.I3(p_s2_o19_4),
.I4(p_s2_o19_5),
.I5(p_s2_o20_0));

/////////STEP3----ORDER20////////////

wire p_s3_o21_1;
wire p_s3_o20_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o20_t198_z0_v0 (
.O6(p_s3_o21_1),
.O5(p_s3_o20_2),
.I0(p_s2_o20_1),
.I1(p_s2_o20_2),
.I2(p_s2_o20_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER21////////////

wire p_s3_o21_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o21_t229_z0_v0 (
.O6(p_s3_o21_2),
.O5(),
.I0(p_s2_o21_0),
.I1(p_s2_o21_1),
.I2(p_s2_o21_2),
.I3(p_s2_o21_3),
.I4(p_s2_o21_4),
.I5(p_s2_o22_0));

wire p_s3_o22_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o21_t229_z1_v0 (
.O6(p_s3_o22_0),
.O5(),
.I0(p_s2_o21_0),
.I1(p_s2_o21_1),
.I2(p_s2_o21_2),
.I3(p_s2_o21_3),
.I4(p_s2_o21_4),
.I5(p_s2_o22_0));

wire p_s3_o23_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o21_t229_z2_v0 (
.O6(p_s3_o23_0),
.O5(),
.I0(p_s2_o21_0),
.I1(p_s2_o21_1),
.I2(p_s2_o21_2),
.I3(p_s2_o21_3),
.I4(p_s2_o21_4),
.I5(p_s2_o22_0));

/////////STEP3----ORDER22////////////

wire p_s3_o22_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o22_t230_z0_v0 (
.O6(p_s3_o22_1),
.O5(),
.I0(p_s2_o22_1),
.I1(p_s2_o22_2),
.I2(p_s2_o22_3),
.I3(p_s2_o22_4),
.I4(p_s2_o22_5),
.I5(p_s2_o23_0));

wire p_s3_o23_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o22_t230_z1_v0 (
.O6(p_s3_o23_1),
.O5(),
.I0(p_s2_o22_1),
.I1(p_s2_o22_2),
.I2(p_s2_o22_3),
.I3(p_s2_o22_4),
.I4(p_s2_o22_5),
.I5(p_s2_o23_0));

wire p_s3_o24_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o22_t230_z2_v0 (
.O6(p_s3_o24_0),
.O5(),
.I0(p_s2_o22_1),
.I1(p_s2_o22_2),
.I2(p_s2_o22_3),
.I3(p_s2_o22_4),
.I4(p_s2_o22_5),
.I5(p_s2_o23_0));

/////////STEP3----ORDER23////////////

wire p_s3_o24_1;
wire p_s3_o23_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o23_t199_z0_v0 (
.O6(p_s3_o24_1),
.O5(p_s3_o23_2),
.I0(p_s2_o23_1),
.I1(p_s2_o23_2),
.I2(p_s2_o23_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER24////////////

wire p_s3_o24_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o24_t231_z0_v0 (
.O6(p_s3_o24_2),
.O5(),
.I0(p_s2_o24_0),
.I1(p_s2_o24_1),
.I2(p_s2_o24_2),
.I3(p_s2_o24_3),
.I4(p_s2_o24_4),
.I5(p_s2_o25_0));

wire p_s3_o25_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o24_t231_z1_v0 (
.O6(p_s3_o25_0),
.O5(),
.I0(p_s2_o24_0),
.I1(p_s2_o24_1),
.I2(p_s2_o24_2),
.I3(p_s2_o24_3),
.I4(p_s2_o24_4),
.I5(p_s2_o25_0));

wire p_s3_o26_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o24_t231_z2_v0 (
.O6(p_s3_o26_0),
.O5(),
.I0(p_s2_o24_0),
.I1(p_s2_o24_1),
.I2(p_s2_o24_2),
.I3(p_s2_o24_3),
.I4(p_s2_o24_4),
.I5(p_s2_o25_0));

/////////STEP3----ORDER25////////////

wire p_s3_o25_1;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s3_o25_t221_z0_v0 (
.O6(p_s3_o25_1),
.O5(),
.I0(p_s2_o25_1),
.I1(p_s2_o25_2),
.I2(p_s2_o25_3),
.I3(p_s2_o25_4),
.I4(p_s2_o25_5),
.I5(p_s0_o25_11));

wire p_s3_o26_1;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s3_o25_t221_z1_v0 (
.O6(p_s3_o26_1),
.O5(),
.I0(p_s2_o25_1),
.I1(p_s2_o25_2),
.I2(p_s2_o25_3),
.I3(p_s2_o25_4),
.I4(p_s2_o25_5),
.I5(p_s0_o25_11));

wire p_s3_o27_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s3_o25_t221_z2_v0 (
.O6(p_s3_o27_0),
.O5(),
.I0(p_s2_o25_1),
.I1(p_s2_o25_2),
.I2(p_s2_o25_3),
.I3(p_s2_o25_4),
.I4(p_s2_o25_5),
.I5(p_s0_o25_11));

/////////STEP3----ORDER26////////////

wire p_s3_o27_1;
wire p_s3_o26_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o26_t200_z0_v0 (
.O6(p_s3_o27_1),
.O5(p_s3_o26_2),
.I0(p_s2_o26_0),
.I1(p_s2_o26_1),
.I2(p_s2_o26_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o27_2;
wire p_s3_o26_3;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o26_t200_z0_v1 (
.O6(p_s3_o27_2),
.O5(p_s3_o26_3),
.I0(p_s2_o26_3),
.I1(p_s2_o26_4),
.I2(p_s2_o26_5),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER27////////////

wire p_s3_o27_3;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s3_o27_t222_z0_v0 (
.O6(p_s3_o27_3),
.O5(),
.I0(p_s2_o27_0),
.I1(p_s2_o27_1),
.I2(p_s2_o27_2),
.I3(p_s2_o27_3),
.I4(p_s2_o27_4),
.I5(p_s2_o27_5));

wire p_s3_o28_0;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s3_o27_t222_z1_v0 (
.O6(p_s3_o28_0),
.O5(),
.I0(p_s2_o27_0),
.I1(p_s2_o27_1),
.I2(p_s2_o27_2),
.I3(p_s2_o27_3),
.I4(p_s2_o27_4),
.I5(p_s2_o27_5));

wire p_s3_o29_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s3_o27_t222_z2_v0 (
.O6(p_s3_o29_0),
.O5(),
.I0(p_s2_o27_0),
.I1(p_s2_o27_1),
.I2(p_s2_o27_2),
.I3(p_s2_o27_3),
.I4(p_s2_o27_4),
.I5(p_s2_o27_5));

/////////STEP3----ORDER28////////////

wire p_s3_o28_1;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s3_o28_t223_z0_v0 (
.O6(p_s3_o28_1),
.O5(),
.I0(p_s2_o28_0),
.I1(p_s2_o28_1),
.I2(p_s2_o28_2),
.I3(p_s2_o28_3),
.I4(p_s2_o28_4),
.I5(p_s2_o28_5));

wire p_s3_o29_1;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s3_o28_t223_z1_v0 (
.O6(p_s3_o29_1),
.O5(),
.I0(p_s2_o28_0),
.I1(p_s2_o28_1),
.I2(p_s2_o28_2),
.I3(p_s2_o28_3),
.I4(p_s2_o28_4),
.I5(p_s2_o28_5));

wire p_s3_o30_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s3_o28_t223_z2_v0 (
.O6(p_s3_o30_0),
.O5(),
.I0(p_s2_o28_0),
.I1(p_s2_o28_1),
.I2(p_s2_o28_2),
.I3(p_s2_o28_3),
.I4(p_s2_o28_4),
.I5(p_s2_o28_5));

/////////STEP3----ORDER29////////////

wire p_s3_o29_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o29_t232_z0_v0 (
.O6(p_s3_o29_2),
.O5(),
.I0(p_s2_o29_0),
.I1(p_s2_o29_1),
.I2(p_s2_o29_2),
.I3(p_s2_o29_3),
.I4(p_s2_o29_4),
.I5(p_s2_o30_0));

wire p_s3_o30_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o29_t232_z1_v0 (
.O6(p_s3_o30_1),
.O5(),
.I0(p_s2_o29_0),
.I1(p_s2_o29_1),
.I2(p_s2_o29_2),
.I3(p_s2_o29_3),
.I4(p_s2_o29_4),
.I5(p_s2_o30_0));

wire p_s3_o31_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o29_t232_z2_v0 (
.O6(p_s3_o31_0),
.O5(),
.I0(p_s2_o29_0),
.I1(p_s2_o29_1),
.I2(p_s2_o29_2),
.I3(p_s2_o29_3),
.I4(p_s2_o29_4),
.I5(p_s2_o30_0));

/////////STEP3----ORDER30////////////

wire p_s3_o30_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o30_t233_z0_v0 (
.O6(p_s3_o30_2),
.O5(),
.I0(p_s2_o30_1),
.I1(p_s2_o30_2),
.I2(p_s2_o30_3),
.I3(p_s2_o30_4),
.I4(p_s2_o30_5),
.I5(p_s2_o31_0));

wire p_s3_o31_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o30_t233_z1_v0 (
.O6(p_s3_o31_1),
.O5(),
.I0(p_s2_o30_1),
.I1(p_s2_o30_2),
.I2(p_s2_o30_3),
.I3(p_s2_o30_4),
.I4(p_s2_o30_5),
.I5(p_s2_o31_0));

wire p_s3_o32_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o30_t233_z2_v0 (
.O6(p_s3_o32_0),
.O5(),
.I0(p_s2_o30_1),
.I1(p_s2_o30_2),
.I2(p_s2_o30_3),
.I3(p_s2_o30_4),
.I4(p_s2_o30_5),
.I5(p_s2_o31_0));

/////////STEP3----ORDER31////////////

wire p_s3_o31_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o31_t234_z0_v0 (
.O6(p_s3_o31_2),
.O5(),
.I0(p_s2_o31_1),
.I1(p_s2_o31_2),
.I2(p_s2_o31_3),
.I3(p_s2_o31_4),
.I4(p_s2_o31_5),
.I5(p_s2_o32_0));

wire p_s3_o32_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o31_t234_z1_v0 (
.O6(p_s3_o32_1),
.O5(),
.I0(p_s2_o31_1),
.I1(p_s2_o31_2),
.I2(p_s2_o31_3),
.I3(p_s2_o31_4),
.I4(p_s2_o31_5),
.I5(p_s2_o32_0));

wire p_s3_o33_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o31_t234_z2_v0 (
.O6(p_s3_o33_0),
.O5(),
.I0(p_s2_o31_1),
.I1(p_s2_o31_2),
.I2(p_s2_o31_3),
.I3(p_s2_o31_4),
.I4(p_s2_o31_5),
.I5(p_s2_o32_0));

/////////STEP3----ORDER32////////////

wire p_s3_o32_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o32_t235_z0_v0 (
.O6(p_s3_o32_2),
.O5(),
.I0(p_s2_o32_1),
.I1(p_s2_o32_2),
.I2(p_s2_o32_3),
.I3(p_s2_o32_4),
.I4(p_s2_o32_5),
.I5(p_s2_o33_0));

wire p_s3_o33_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o32_t235_z1_v0 (
.O6(p_s3_o33_1),
.O5(),
.I0(p_s2_o32_1),
.I1(p_s2_o32_2),
.I2(p_s2_o32_3),
.I3(p_s2_o32_4),
.I4(p_s2_o32_5),
.I5(p_s2_o33_0));

wire p_s3_o34_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o32_t235_z2_v0 (
.O6(p_s3_o34_0),
.O5(),
.I0(p_s2_o32_1),
.I1(p_s2_o32_2),
.I2(p_s2_o32_3),
.I3(p_s2_o32_4),
.I4(p_s2_o32_5),
.I5(p_s2_o33_0));

/////////STEP3----ORDER33////////////

wire p_s3_o34_1;
wire p_s3_o33_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o33_t201_z0_v0 (
.O6(p_s3_o34_1),
.O5(p_s3_o33_2),
.I0(p_s2_o33_1),
.I1(p_s2_o33_2),
.I2(p_s2_o33_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER34////////////

wire p_s3_o34_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o34_t236_z0_v0 (
.O6(p_s3_o34_2),
.O5(),
.I0(p_s2_o34_0),
.I1(p_s2_o34_1),
.I2(p_s2_o34_2),
.I3(p_s2_o34_3),
.I4(p_s2_o34_4),
.I5(p_s2_o35_0));

wire p_s3_o35_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o34_t236_z1_v0 (
.O6(p_s3_o35_0),
.O5(),
.I0(p_s2_o34_0),
.I1(p_s2_o34_1),
.I2(p_s2_o34_2),
.I3(p_s2_o34_3),
.I4(p_s2_o34_4),
.I5(p_s2_o35_0));

wire p_s3_o36_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o34_t236_z2_v0 (
.O6(p_s3_o36_0),
.O5(),
.I0(p_s2_o34_0),
.I1(p_s2_o34_1),
.I2(p_s2_o34_2),
.I3(p_s2_o34_3),
.I4(p_s2_o34_4),
.I5(p_s2_o35_0));

/////////STEP3----ORDER35////////////

wire p_s3_o35_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o35_t237_z0_v0 (
.O6(p_s3_o35_1),
.O5(),
.I0(p_s2_o35_1),
.I1(p_s2_o35_2),
.I2(p_s2_o35_3),
.I3(p_s2_o35_4),
.I4(p_s2_o35_5),
.I5(p_s2_o36_0));

wire p_s3_o36_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o35_t237_z1_v0 (
.O6(p_s3_o36_1),
.O5(),
.I0(p_s2_o35_1),
.I1(p_s2_o35_2),
.I2(p_s2_o35_3),
.I3(p_s2_o35_4),
.I4(p_s2_o35_5),
.I5(p_s2_o36_0));

wire p_s3_o37_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o35_t237_z2_v0 (
.O6(p_s3_o37_0),
.O5(),
.I0(p_s2_o35_1),
.I1(p_s2_o35_2),
.I2(p_s2_o35_3),
.I3(p_s2_o35_4),
.I4(p_s2_o35_5),
.I5(p_s2_o36_0));

/////////STEP3----ORDER36////////////

wire p_s3_o36_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o36_t238_z0_v0 (
.O6(p_s3_o36_2),
.O5(),
.I0(p_s2_o36_1),
.I1(p_s2_o36_2),
.I2(p_s2_o36_3),
.I3(p_s2_o36_4),
.I4(p_s2_o36_5),
.I5(p_s2_o37_0));

wire p_s3_o37_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o36_t238_z1_v0 (
.O6(p_s3_o37_1),
.O5(),
.I0(p_s2_o36_1),
.I1(p_s2_o36_2),
.I2(p_s2_o36_3),
.I3(p_s2_o36_4),
.I4(p_s2_o36_5),
.I5(p_s2_o37_0));

wire p_s3_o38_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o36_t238_z2_v0 (
.O6(p_s3_o38_0),
.O5(),
.I0(p_s2_o36_1),
.I1(p_s2_o36_2),
.I2(p_s2_o36_3),
.I3(p_s2_o36_4),
.I4(p_s2_o36_5),
.I5(p_s2_o37_0));

/////////STEP3----ORDER37////////////

wire p_s3_o37_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o37_t239_z0_v0 (
.O6(p_s3_o37_2),
.O5(),
.I0(p_s2_o37_1),
.I1(p_s2_o37_2),
.I2(p_s2_o37_3),
.I3(p_s2_o37_4),
.I4(p_s2_o37_5),
.I5(p_s2_o38_0));

wire p_s3_o38_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o37_t239_z1_v0 (
.O6(p_s3_o38_1),
.O5(),
.I0(p_s2_o37_1),
.I1(p_s2_o37_2),
.I2(p_s2_o37_3),
.I3(p_s2_o37_4),
.I4(p_s2_o37_5),
.I5(p_s2_o38_0));

wire p_s3_o39_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o37_t239_z2_v0 (
.O6(p_s3_o39_0),
.O5(),
.I0(p_s2_o37_1),
.I1(p_s2_o37_2),
.I2(p_s2_o37_3),
.I3(p_s2_o37_4),
.I4(p_s2_o37_5),
.I5(p_s2_o38_0));

/////////STEP3----ORDER38////////////

wire p_s3_o38_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o38_t240_z0_v0 (
.O6(p_s3_o38_2),
.O5(),
.I0(p_s2_o38_1),
.I1(p_s2_o38_2),
.I2(p_s2_o38_3),
.I3(p_s2_o38_4),
.I4(p_s2_o38_5),
.I5(p_s2_o39_0));

wire p_s3_o39_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o38_t240_z1_v0 (
.O6(p_s3_o39_1),
.O5(),
.I0(p_s2_o38_1),
.I1(p_s2_o38_2),
.I2(p_s2_o38_3),
.I3(p_s2_o38_4),
.I4(p_s2_o38_5),
.I5(p_s2_o39_0));

wire p_s3_o40_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o38_t240_z2_v0 (
.O6(p_s3_o40_0),
.O5(),
.I0(p_s2_o38_1),
.I1(p_s2_o38_2),
.I2(p_s2_o38_3),
.I3(p_s2_o38_4),
.I4(p_s2_o38_5),
.I5(p_s2_o39_0));

/////////STEP3----ORDER39////////////

wire p_s3_o40_1;
wire p_s3_o39_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o39_t202_z0_v0 (
.O6(p_s3_o40_1),
.O5(p_s3_o39_2),
.I0(p_s2_o39_1),
.I1(p_s2_o39_2),
.I2(p_s2_o39_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER40////////////

wire p_s3_o40_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o40_t241_z0_v0 (
.O6(p_s3_o40_2),
.O5(),
.I0(p_s2_o40_0),
.I1(p_s2_o40_1),
.I2(p_s2_o40_2),
.I3(p_s2_o40_3),
.I4(p_s2_o40_4),
.I5(p_s2_o41_0));

wire p_s3_o41_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o40_t241_z1_v0 (
.O6(p_s3_o41_0),
.O5(),
.I0(p_s2_o40_0),
.I1(p_s2_o40_1),
.I2(p_s2_o40_2),
.I3(p_s2_o40_3),
.I4(p_s2_o40_4),
.I5(p_s2_o41_0));

wire p_s3_o42_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o40_t241_z2_v0 (
.O6(p_s3_o42_0),
.O5(),
.I0(p_s2_o40_0),
.I1(p_s2_o40_1),
.I2(p_s2_o40_2),
.I3(p_s2_o40_3),
.I4(p_s2_o40_4),
.I5(p_s2_o41_0));

/////////STEP3----ORDER41////////////

wire p_s3_o41_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o41_t242_z0_v0 (
.O6(p_s3_o41_1),
.O5(),
.I0(p_s2_o41_1),
.I1(p_s2_o41_2),
.I2(p_s2_o41_3),
.I3(p_s2_o41_4),
.I4(p_s2_o41_5),
.I5(p_s2_o42_0));

wire p_s3_o42_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o41_t242_z1_v0 (
.O6(p_s3_o42_1),
.O5(),
.I0(p_s2_o41_1),
.I1(p_s2_o41_2),
.I2(p_s2_o41_3),
.I3(p_s2_o41_4),
.I4(p_s2_o41_5),
.I5(p_s2_o42_0));

wire p_s3_o43_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o41_t242_z2_v0 (
.O6(p_s3_o43_0),
.O5(),
.I0(p_s2_o41_1),
.I1(p_s2_o41_2),
.I2(p_s2_o41_3),
.I3(p_s2_o41_4),
.I4(p_s2_o41_5),
.I5(p_s2_o42_0));

/////////STEP3----ORDER42////////////

wire p_s3_o43_1;
wire p_s3_o42_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o42_t203_z0_v0 (
.O6(p_s3_o43_1),
.O5(p_s3_o42_2),
.I0(p_s2_o42_1),
.I1(p_s2_o42_2),
.I2(p_s2_o42_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER43////////////

wire p_s3_o43_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o43_t243_z0_v0 (
.O6(p_s3_o43_2),
.O5(),
.I0(p_s2_o43_0),
.I1(p_s2_o43_1),
.I2(p_s2_o43_2),
.I3(p_s2_o43_3),
.I4(p_s2_o43_4),
.I5(p_s2_o44_0));

wire p_s3_o44_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o43_t243_z1_v0 (
.O6(p_s3_o44_0),
.O5(),
.I0(p_s2_o43_0),
.I1(p_s2_o43_1),
.I2(p_s2_o43_2),
.I3(p_s2_o43_3),
.I4(p_s2_o43_4),
.I5(p_s2_o44_0));

wire p_s3_o45_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o43_t243_z2_v0 (
.O6(p_s3_o45_0),
.O5(),
.I0(p_s2_o43_0),
.I1(p_s2_o43_1),
.I2(p_s2_o43_2),
.I3(p_s2_o43_3),
.I4(p_s2_o43_4),
.I5(p_s2_o44_0));

/////////STEP3----ORDER44////////////

wire p_s3_o44_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o44_t244_z0_v0 (
.O6(p_s3_o44_1),
.O5(),
.I0(p_s2_o44_1),
.I1(p_s2_o44_2),
.I2(p_s2_o44_3),
.I3(p_s2_o44_4),
.I4(p_s2_o44_5),
.I5(p_s2_o45_0));

wire p_s3_o45_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o44_t244_z1_v0 (
.O6(p_s3_o45_1),
.O5(),
.I0(p_s2_o44_1),
.I1(p_s2_o44_2),
.I2(p_s2_o44_3),
.I3(p_s2_o44_4),
.I4(p_s2_o44_5),
.I5(p_s2_o45_0));

wire p_s3_o46_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o44_t244_z2_v0 (
.O6(p_s3_o46_0),
.O5(),
.I0(p_s2_o44_1),
.I1(p_s2_o44_2),
.I2(p_s2_o44_3),
.I3(p_s2_o44_4),
.I4(p_s2_o44_5),
.I5(p_s2_o45_0));

/////////STEP3----ORDER45////////////

wire p_s3_o45_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o45_t245_z0_v0 (
.O6(p_s3_o45_2),
.O5(),
.I0(p_s2_o45_1),
.I1(p_s2_o45_2),
.I2(p_s2_o45_3),
.I3(p_s2_o45_4),
.I4(p_s2_o45_5),
.I5(p_s2_o46_0));

wire p_s3_o46_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o45_t245_z1_v0 (
.O6(p_s3_o46_1),
.O5(),
.I0(p_s2_o45_1),
.I1(p_s2_o45_2),
.I2(p_s2_o45_3),
.I3(p_s2_o45_4),
.I4(p_s2_o45_5),
.I5(p_s2_o46_0));

wire p_s3_o47_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o45_t245_z2_v0 (
.O6(p_s3_o47_0),
.O5(),
.I0(p_s2_o45_1),
.I1(p_s2_o45_2),
.I2(p_s2_o45_3),
.I3(p_s2_o45_4),
.I4(p_s2_o45_5),
.I5(p_s2_o46_0));

/////////STEP3----ORDER46////////////

wire p_s3_o46_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o46_t246_z0_v0 (
.O6(p_s3_o46_2),
.O5(),
.I0(p_s2_o46_1),
.I1(p_s2_o46_2),
.I2(p_s2_o46_3),
.I3(p_s2_o46_4),
.I4(p_s2_o46_5),
.I5(p_s2_o47_0));

wire p_s3_o47_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o46_t246_z1_v0 (
.O6(p_s3_o47_1),
.O5(),
.I0(p_s2_o46_1),
.I1(p_s2_o46_2),
.I2(p_s2_o46_3),
.I3(p_s2_o46_4),
.I4(p_s2_o46_5),
.I5(p_s2_o47_0));

wire p_s3_o48_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o46_t246_z2_v0 (
.O6(p_s3_o48_0),
.O5(),
.I0(p_s2_o46_1),
.I1(p_s2_o46_2),
.I2(p_s2_o46_3),
.I3(p_s2_o46_4),
.I4(p_s2_o46_5),
.I5(p_s2_o47_0));

/////////STEP3----ORDER47////////////

wire p_s3_o48_1;
wire p_s3_o47_2;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o47_t208_z0_v0 (
.O6(p_s3_o48_1),
.O5(p_s3_o47_2),
.I0(a[20]),
.I1(b[30]),
.I2(p_s2_o47_1),
.I3(p_s2_o47_2),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o48_2;
wire p_s3_o47_3;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o47_t208_z0_v1 (
.O6(p_s3_o48_2),
.O5(p_s3_o47_3),
.I0(a[19]),
.I1(b[31]),
.I2(p_s2_o47_3),
.I3(p_s2_o47_4),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER48////////////

wire p_s3_o48_3;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o48_t247_z0_v0 (
.O6(p_s3_o48_3),
.O5(),
.I0(p_s2_o48_0),
.I1(p_s2_o48_1),
.I2(p_s2_o48_2),
.I3(p_s2_o48_3),
.I4(p_s1_o48_5),
.I5(p_s2_o49_0));

wire p_s3_o49_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o48_t247_z1_v0 (
.O6(p_s3_o49_0),
.O5(),
.I0(p_s2_o48_0),
.I1(p_s2_o48_1),
.I2(p_s2_o48_2),
.I3(p_s2_o48_3),
.I4(p_s1_o48_5),
.I5(p_s2_o49_0));

wire p_s3_o50_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o48_t247_z2_v0 (
.O6(p_s3_o50_0),
.O5(),
.I0(p_s2_o48_0),
.I1(p_s2_o48_1),
.I2(p_s2_o48_2),
.I3(p_s2_o48_3),
.I4(p_s1_o48_5),
.I5(p_s2_o49_0));

/////////STEP3----ORDER49////////////

wire p_s3_o49_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o49_t248_z0_v0 (
.O6(p_s3_o49_1),
.O5(),
.I0(p_s2_o49_1),
.I1(p_s2_o49_2),
.I2(p_s2_o49_3),
.I3(p_s2_o49_4),
.I4(p_s2_o49_5),
.I5(p_s2_o50_0));

wire p_s3_o50_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o49_t248_z1_v0 (
.O6(p_s3_o50_1),
.O5(),
.I0(p_s2_o49_1),
.I1(p_s2_o49_2),
.I2(p_s2_o49_3),
.I3(p_s2_o49_4),
.I4(p_s2_o49_5),
.I5(p_s2_o50_0));

wire p_s3_o51_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o49_t248_z2_v0 (
.O6(p_s3_o51_0),
.O5(),
.I0(p_s2_o49_1),
.I1(p_s2_o49_2),
.I2(p_s2_o49_3),
.I3(p_s2_o49_4),
.I4(p_s2_o49_5),
.I5(p_s2_o50_0));

/////////STEP3----ORDER50////////////

wire p_s3_o51_1;
wire p_s3_o50_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o50_t204_z0_v0 (
.O6(p_s3_o51_1),
.O5(p_s3_o50_2),
.I0(p_s2_o50_1),
.I1(p_s2_o50_2),
.I2(p_s2_o50_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o51_2;
wire p_s3_o50_3;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o50_t209_z0_v0 (
.O6(p_s3_o51_2),
.O5(p_s3_o50_3),
.I0(a[22]),
.I1(b[31]),
.I2(p_s2_o50_4),
.I3(p_s2_o50_5),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER51////////////

wire p_s3_o51_3;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o51_t249_z0_v0 (
.O6(p_s3_o51_3),
.O5(),
.I0(p_s2_o51_0),
.I1(p_s2_o51_1),
.I2(p_s2_o51_2),
.I3(p_s2_o51_3),
.I4(p_s1_o51_1),
.I5(p_s2_o52_0));

wire p_s3_o52_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o51_t249_z1_v0 (
.O6(p_s3_o52_0),
.O5(),
.I0(p_s2_o51_0),
.I1(p_s2_o51_1),
.I2(p_s2_o51_2),
.I3(p_s2_o51_3),
.I4(p_s1_o51_1),
.I5(p_s2_o52_0));

wire p_s3_o53_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o51_t249_z2_v0 (
.O6(p_s3_o53_0),
.O5(),
.I0(p_s2_o51_0),
.I1(p_s2_o51_1),
.I2(p_s2_o51_2),
.I3(p_s2_o51_3),
.I4(p_s1_o51_1),
.I5(p_s2_o52_0));

/////////STEP3----ORDER52////////////

wire p_s3_o53_1;
wire p_s3_o52_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o52_t205_z0_v0 (
.O6(p_s3_o53_1),
.O5(p_s3_o52_1),
.I0(p_s2_o52_1),
.I1(p_s2_o52_2),
.I2(p_s2_o52_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER53////////////

wire p_s3_o54_0;
wire p_s3_o53_2;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o53_t210_z0_v0 (
.O6(p_s3_o54_0),
.O5(p_s3_o53_2),
.I0(a[29]),
.I1(b[27]),
.I2(p_s2_o53_0),
.I3(p_s2_o53_1),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o54_1;
wire p_s3_o53_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o53_t216_z0_v0 (
.O6(p_s3_o54_1),
.O5(p_s3_o53_3),
.I0(a[28]),
.I1(b[28]),
.I2(a[27]),
.I3(b[29]),
.I4(p_s2_o53_2),
.I5(1'b1));

wire p_s3_o54_2;
wire p_s3_o53_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o53_t216_z0_v1 (
.O6(p_s3_o54_2),
.O5(p_s3_o53_4),
.I0(a[26]),
.I1(b[30]),
.I2(a[25]),
.I3(b[31]),
.I4(p_s2_o53_3),
.I5(1'b1));

/////////STEP3----ORDER54////////////

wire p_s3_o55_0;
wire p_s3_o54_3;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o54_t211_z0_v0 (
.O6(p_s3_o55_0),
.O5(p_s3_o54_3),
.I0(a[26]),
.I1(b[31]),
.I2(p_s2_o54_0),
.I3(p_s1_o54_0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER55////////////

wire p_s3_o56_0;
wire p_s3_o55_1;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o55_t212_z0_v0 (
.O6(p_s3_o56_0),
.O5(p_s3_o55_1),
.I0(a[27]),
.I1(b[31]),
.I2(p_s2_o55_0),
.I3(p_s1_o55_1),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER56////////////

wire p_s3_o57_0;
wire p_s3_o56_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o56_t217_z0_v0 (
.O6(p_s3_o57_0),
.O5(p_s3_o56_1),
.I0(a[29]),
.I1(b[30]),
.I2(a[28]),
.I3(b[31]),
.I4(p_s2_o56_0),
.I5(1'b1));

/////////STEP3----ORDER57////////////

wire p_s3_o58_0;
wire p_s3_o57_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o57_t218_z0_v0 (
.O6(p_s3_o58_0),
.O5(p_s3_o57_1),
.I0(a[31]),
.I1(b[29]),
.I2(a[30]),
.I3(b[30]),
.I4(p_s2_o57_0),
.I5(1'b1));

/////////STEP3----ORDER58////////////

/////////STEP3----ORDER59////////////

/////////STEP4----ORDER0////////////

LUT6_2 #(
.INIT(64'h8778877808800880)
) LUT6_2_inst_oo0 (
.O6(P[0]),
.O5(G[0]),
.I0(a[0]),
.I1(b[3]),
.I2(C0),
.I3(p_s0_o0_0),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER1////////////

LUT6_2 #(
.INIT(64'h8778787878000000)
) LUT6_2_inst_oo1 (
.O6(P[1]),
.O5(G[1]),
.I0(a[0]),
.I1(b[4]),
.I2(p_s2_o1_0),
.I3(C0),
.I4(p_s0_o0_0),
.I5(1'b1));

/////////STEP4----ORDER2////////////

LUT6_2 #(
.INIT(64'h9666666660000000)
) LUT6_2_inst_oo2 (
.O6(P[2]),
.O5(G[2]),
.I0(p_s3_o2_0),
.I1(p_s3_o2_1),
.I2(a[0]),
.I3(b[4]),
.I4(p_s2_o1_0),
.I5(1'b1));

/////////STEP4----ORDER3////////////

wire p_s4_o4_0;
wire p_s4_o3_0;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s4_o3_t250_z0_v0 (
.O6(p_s4_o4_0),
.O5(p_s4_o3_0),
.I0(p_s3_o3_0),
.I1(p_s3_o3_1),
.I2(p_s2_o3_0),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo3 (
.O6(P[3]),
.O5(G[3]),
.I0(p_s4_o3_0),
.I1(p_s2_o3_1),
.I2(p_s3_o2_0),
.I3(p_s3_o2_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER4////////////

wire p_s4_o5_0;
wire p_s4_o4_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o4_t271_z0_v0 (
.O6(p_s4_o5_0),
.O5(p_s4_o4_1),
.I0(p_s3_o4_0),
.I1(p_s1_o4_1),
.I2(p_s1_o4_2),
.I3(p_s3_o5_0),
.I4(p_s3_o5_1),
.I5(1'b1));

wire p_s4_o6_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o4_t271_z1_v0 (
.O6(p_s4_o6_0),
.O5(),
.I0(p_s3_o4_0),
.I1(p_s1_o4_1),
.I2(p_s1_o4_2),
.I3(p_s3_o5_0),
.I4(p_s3_o5_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo4 (
.O6(P[4]),
.O5(G[4]),
.I0(p_s4_o4_0),
.I1(p_s4_o4_1),
.I2(p_s4_o3_0),
.I3(p_s2_o3_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER5////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo5 (
.O6(P[5]),
.O5(G[5]),
.I0(p_s4_o5_0),
.I1(p_s2_o5_2),
.I2(p_s4_o4_0),
.I3(p_s4_o4_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER6////////////

wire p_s4_o6_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o6_t256_z0_v0 (
.O6(p_s4_o6_1),
.O5(),
.I0(p_s3_o6_0),
.I1(p_s3_o6_1),
.I2(p_s3_o6_2),
.I3(p_s3_o6_3),
.I4(p_s3_o6_4),
.I5(p_s3_o7_0));

wire p_s4_o7_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o6_t256_z1_v0 (
.O6(p_s4_o7_0),
.O5(),
.I0(p_s3_o6_0),
.I1(p_s3_o6_1),
.I2(p_s3_o6_2),
.I3(p_s3_o6_3),
.I4(p_s3_o6_4),
.I5(p_s3_o7_0));

wire p_s4_o8_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o6_t256_z2_v0 (
.O6(p_s4_o8_0),
.O5(),
.I0(p_s3_o6_0),
.I1(p_s3_o6_1),
.I2(p_s3_o6_2),
.I3(p_s3_o6_3),
.I4(p_s3_o6_4),
.I5(p_s3_o7_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo6 (
.O6(P[6]),
.O5(G[6]),
.I0(p_s4_o6_0),
.I1(p_s4_o6_1),
.I2(p_s4_o5_0),
.I3(p_s2_o5_2),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER7////////////

wire p_s4_o7_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o7_t257_z0_v0 (
.O6(p_s4_o7_1),
.O5(),
.I0(p_s3_o7_1),
.I1(p_s3_o7_2),
.I2(p_s3_o7_3),
.I3(p_s2_o7_0),
.I4(p_s2_o7_1),
.I5(p_s3_o8_0));

wire p_s4_o8_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o7_t257_z1_v0 (
.O6(p_s4_o8_1),
.O5(),
.I0(p_s3_o7_1),
.I1(p_s3_o7_2),
.I2(p_s3_o7_3),
.I3(p_s2_o7_0),
.I4(p_s2_o7_1),
.I5(p_s3_o8_0));

wire p_s4_o9_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o7_t257_z2_v0 (
.O6(p_s4_o9_0),
.O5(),
.I0(p_s3_o7_1),
.I1(p_s3_o7_2),
.I2(p_s3_o7_3),
.I3(p_s2_o7_0),
.I4(p_s2_o7_1),
.I5(p_s3_o8_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo7 (
.O6(P[7]),
.O5(G[7]),
.I0(p_s4_o7_0),
.I1(p_s4_o7_1),
.I2(p_s4_o6_0),
.I3(p_s4_o6_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER8////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo8 (
.O6(P[8]),
.O5(G[8]),
.I0(p_s4_o8_0),
.I1(p_s4_o8_1),
.I2(p_s4_o7_0),
.I3(p_s4_o7_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER9////////////

wire p_s4_o9_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o9_t258_z0_v0 (
.O6(p_s4_o9_1),
.O5(),
.I0(p_s3_o9_0),
.I1(p_s3_o9_1),
.I2(p_s3_o9_2),
.I3(p_s2_o9_5),
.I4(p_s2_o9_6),
.I5(p_s3_o10_0));

wire p_s4_o10_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o9_t258_z1_v0 (
.O6(p_s4_o10_0),
.O5(),
.I0(p_s3_o9_0),
.I1(p_s3_o9_1),
.I2(p_s3_o9_2),
.I3(p_s2_o9_5),
.I4(p_s2_o9_6),
.I5(p_s3_o10_0));

wire p_s4_o11_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o9_t258_z2_v0 (
.O6(p_s4_o11_0),
.O5(),
.I0(p_s3_o9_0),
.I1(p_s3_o9_1),
.I2(p_s3_o9_2),
.I3(p_s2_o9_5),
.I4(p_s2_o9_6),
.I5(p_s3_o10_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo9 (
.O6(P[9]),
.O5(G[9]),
.I0(p_s4_o9_0),
.I1(p_s4_o9_1),
.I2(p_s4_o8_0),
.I3(p_s4_o8_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER10////////////

wire p_s4_o11_1;
wire p_s4_o10_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o10_t272_z0_v0 (
.O6(p_s4_o11_1),
.O5(p_s4_o10_1),
.I0(p_s3_o10_1),
.I1(p_s3_o10_2),
.I2(p_s3_o10_3),
.I3(p_s3_o11_0),
.I4(p_s3_o11_1),
.I5(1'b1));

wire p_s4_o12_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o10_t272_z1_v0 (
.O6(p_s4_o12_0),
.O5(),
.I0(p_s3_o10_1),
.I1(p_s3_o10_2),
.I2(p_s3_o10_3),
.I3(p_s3_o11_0),
.I4(p_s3_o11_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo10 (
.O6(P[10]),
.O5(G[10]),
.I0(p_s4_o10_0),
.I1(p_s4_o10_1),
.I2(p_s4_o9_0),
.I3(p_s4_o9_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER11////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo11 (
.O6(P[11]),
.O5(G[11]),
.I0(p_s4_o11_0),
.I1(p_s4_o11_1),
.I2(p_s4_o10_0),
.I3(p_s4_o10_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER12////////////

wire p_s4_o12_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o12_t259_z0_v0 (
.O6(p_s4_o12_1),
.O5(),
.I0(p_s3_o12_0),
.I1(p_s3_o12_1),
.I2(p_s3_o12_2),
.I3(p_s2_o12_5),
.I4(p_s2_o12_6),
.I5(p_s3_o13_0));

wire p_s4_o13_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o12_t259_z1_v0 (
.O6(p_s4_o13_0),
.O5(),
.I0(p_s3_o12_0),
.I1(p_s3_o12_1),
.I2(p_s3_o12_2),
.I3(p_s2_o12_5),
.I4(p_s2_o12_6),
.I5(p_s3_o13_0));

wire p_s4_o14_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o12_t259_z2_v0 (
.O6(p_s4_o14_0),
.O5(),
.I0(p_s3_o12_0),
.I1(p_s3_o12_1),
.I2(p_s3_o12_2),
.I3(p_s2_o12_5),
.I4(p_s2_o12_6),
.I5(p_s3_o13_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo12 (
.O6(P[12]),
.O5(G[12]),
.I0(p_s4_o12_0),
.I1(p_s4_o12_1),
.I2(p_s4_o11_0),
.I3(p_s4_o11_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER13////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo13 (
.O6(P[13]),
.O5(G[13]),
.I0(p_s4_o13_0),
.I1(p_s3_o13_1),
.I2(p_s4_o12_0),
.I3(p_s4_o12_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER14////////////

wire p_s4_o14_1;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s4_o14_t255_z0_v0 (
.O6(p_s4_o14_1),
.O5(),
.I0(p_s3_o14_0),
.I1(p_s3_o14_1),
.I2(p_s2_o14_0),
.I3(p_s2_o14_1),
.I4(p_s1_o14_7),
.I5(p_s0_o14_6));

wire p_s4_o15_0;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s4_o14_t255_z1_v0 (
.O6(p_s4_o15_0),
.O5(),
.I0(p_s3_o14_0),
.I1(p_s3_o14_1),
.I2(p_s2_o14_0),
.I3(p_s2_o14_1),
.I4(p_s1_o14_7),
.I5(p_s0_o14_6));

wire p_s4_o16_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s4_o14_t255_z2_v0 (
.O6(p_s4_o16_0),
.O5(),
.I0(p_s3_o14_0),
.I1(p_s3_o14_1),
.I2(p_s2_o14_0),
.I3(p_s2_o14_1),
.I4(p_s1_o14_7),
.I5(p_s0_o14_6));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo14 (
.O6(P[14]),
.O5(G[14]),
.I0(p_s4_o14_0),
.I1(p_s4_o14_1),
.I2(p_s4_o13_0),
.I3(p_s3_o13_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER15////////////

wire p_s4_o15_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o15_t260_z0_v0 (
.O6(p_s4_o15_1),
.O5(),
.I0(p_s3_o15_0),
.I1(p_s2_o15_0),
.I2(p_s2_o15_1),
.I3(p_s2_o15_2),
.I4(p_s2_o15_3),
.I5(p_s3_o16_0));

wire p_s4_o16_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o15_t260_z1_v0 (
.O6(p_s4_o16_1),
.O5(),
.I0(p_s3_o15_0),
.I1(p_s2_o15_0),
.I2(p_s2_o15_1),
.I3(p_s2_o15_2),
.I4(p_s2_o15_3),
.I5(p_s3_o16_0));

wire p_s4_o17_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o15_t260_z2_v0 (
.O6(p_s4_o17_0),
.O5(),
.I0(p_s3_o15_0),
.I1(p_s2_o15_0),
.I2(p_s2_o15_1),
.I3(p_s2_o15_2),
.I4(p_s2_o15_3),
.I5(p_s3_o16_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo15 (
.O6(P[15]),
.O5(G[15]),
.I0(p_s4_o15_0),
.I1(p_s4_o15_1),
.I2(p_s4_o14_0),
.I3(p_s4_o14_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER16////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo16 (
.O6(P[16]),
.O5(G[16]),
.I0(p_s4_o16_0),
.I1(p_s4_o16_1),
.I2(p_s4_o15_0),
.I3(p_s4_o15_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER17////////////

wire p_s4_o17_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o17_t261_z0_v0 (
.O6(p_s4_o17_1),
.O5(),
.I0(p_s3_o17_0),
.I1(p_s3_o17_1),
.I2(p_s3_o17_2),
.I3(p_s2_o17_6),
.I4(p_s1_o17_10),
.I5(p_s3_o18_0));

wire p_s4_o18_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o17_t261_z1_v0 (
.O6(p_s4_o18_0),
.O5(),
.I0(p_s3_o17_0),
.I1(p_s3_o17_1),
.I2(p_s3_o17_2),
.I3(p_s2_o17_6),
.I4(p_s1_o17_10),
.I5(p_s3_o18_0));

wire p_s4_o19_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o17_t261_z2_v0 (
.O6(p_s4_o19_0),
.O5(),
.I0(p_s3_o17_0),
.I1(p_s3_o17_1),
.I2(p_s3_o17_2),
.I3(p_s2_o17_6),
.I4(p_s1_o17_10),
.I5(p_s3_o18_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo17 (
.O6(P[17]),
.O5(G[17]),
.I0(p_s4_o17_0),
.I1(p_s4_o17_1),
.I2(p_s4_o16_0),
.I3(p_s4_o16_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER18////////////

wire p_s4_o19_1;
wire p_s4_o18_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o18_t273_z0_v0 (
.O6(p_s4_o19_1),
.O5(p_s4_o18_1),
.I0(p_s3_o18_1),
.I1(p_s3_o18_2),
.I2(p_s3_o18_3),
.I3(p_s3_o19_0),
.I4(p_s3_o19_1),
.I5(1'b1));

wire p_s4_o20_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o18_t273_z1_v0 (
.O6(p_s4_o20_0),
.O5(),
.I0(p_s3_o18_1),
.I1(p_s3_o18_2),
.I2(p_s3_o18_3),
.I3(p_s3_o19_0),
.I4(p_s3_o19_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo18 (
.O6(P[18]),
.O5(G[18]),
.I0(p_s4_o18_0),
.I1(p_s4_o18_1),
.I2(p_s4_o17_0),
.I3(p_s4_o17_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER19////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo19 (
.O6(P[19]),
.O5(G[19]),
.I0(p_s4_o19_0),
.I1(p_s4_o19_1),
.I2(p_s4_o18_0),
.I3(p_s4_o18_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER20////////////

wire p_s4_o20_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o20_t262_z0_v0 (
.O6(p_s4_o20_1),
.O5(),
.I0(p_s3_o20_0),
.I1(p_s3_o20_1),
.I2(p_s3_o20_2),
.I3(p_s2_o20_4),
.I4(p_s2_o20_5),
.I5(p_s3_o21_0));

wire p_s4_o21_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o20_t262_z1_v0 (
.O6(p_s4_o21_0),
.O5(),
.I0(p_s3_o20_0),
.I1(p_s3_o20_1),
.I2(p_s3_o20_2),
.I3(p_s2_o20_4),
.I4(p_s2_o20_5),
.I5(p_s3_o21_0));

wire p_s4_o22_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o20_t262_z2_v0 (
.O6(p_s4_o22_0),
.O5(),
.I0(p_s3_o20_0),
.I1(p_s3_o20_1),
.I2(p_s3_o20_2),
.I3(p_s2_o20_4),
.I4(p_s2_o20_5),
.I5(p_s3_o21_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo20 (
.O6(P[20]),
.O5(G[20]),
.I0(p_s4_o20_0),
.I1(p_s4_o20_1),
.I2(p_s4_o19_0),
.I3(p_s4_o19_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER21////////////

wire p_s4_o22_1;
wire p_s4_o21_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o21_t274_z0_v0 (
.O6(p_s4_o22_1),
.O5(p_s4_o21_1),
.I0(p_s3_o21_1),
.I1(p_s3_o21_2),
.I2(p_s2_o21_5),
.I3(p_s3_o22_0),
.I4(p_s3_o22_1),
.I5(1'b1));

wire p_s4_o23_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o21_t274_z1_v0 (
.O6(p_s4_o23_0),
.O5(),
.I0(p_s3_o21_1),
.I1(p_s3_o21_2),
.I2(p_s2_o21_5),
.I3(p_s3_o22_0),
.I4(p_s3_o22_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo21 (
.O6(P[21]),
.O5(G[21]),
.I0(p_s4_o21_0),
.I1(p_s4_o21_1),
.I2(p_s4_o20_0),
.I3(p_s4_o20_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER22////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo22 (
.O6(P[22]),
.O5(G[22]),
.I0(p_s4_o22_0),
.I1(p_s4_o22_1),
.I2(p_s4_o21_0),
.I3(p_s4_o21_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER23////////////

wire p_s4_o23_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o23_t263_z0_v0 (
.O6(p_s4_o23_1),
.O5(),
.I0(p_s3_o23_0),
.I1(p_s3_o23_1),
.I2(p_s3_o23_2),
.I3(p_s2_o23_4),
.I4(p_s2_o23_5),
.I5(p_s3_o24_0));

wire p_s4_o24_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o23_t263_z1_v0 (
.O6(p_s4_o24_0),
.O5(),
.I0(p_s3_o23_0),
.I1(p_s3_o23_1),
.I2(p_s3_o23_2),
.I3(p_s2_o23_4),
.I4(p_s2_o23_5),
.I5(p_s3_o24_0));

wire p_s4_o25_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o23_t263_z2_v0 (
.O6(p_s4_o25_0),
.O5(),
.I0(p_s3_o23_0),
.I1(p_s3_o23_1),
.I2(p_s3_o23_2),
.I3(p_s2_o23_4),
.I4(p_s2_o23_5),
.I5(p_s3_o24_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo23 (
.O6(P[23]),
.O5(G[23]),
.I0(p_s4_o23_0),
.I1(p_s4_o23_1),
.I2(p_s4_o22_0),
.I3(p_s4_o22_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER24////////////

wire p_s4_o25_1;
wire p_s4_o24_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o24_t275_z0_v0 (
.O6(p_s4_o25_1),
.O5(p_s4_o24_1),
.I0(p_s3_o24_1),
.I1(p_s3_o24_2),
.I2(p_s2_o24_5),
.I3(p_s3_o25_0),
.I4(p_s3_o25_1),
.I5(1'b1));

wire p_s4_o26_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o24_t275_z1_v0 (
.O6(p_s4_o26_0),
.O5(),
.I0(p_s3_o24_1),
.I1(p_s3_o24_2),
.I2(p_s2_o24_5),
.I3(p_s3_o25_0),
.I4(p_s3_o25_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo24 (
.O6(P[24]),
.O5(G[24]),
.I0(p_s4_o24_0),
.I1(p_s4_o24_1),
.I2(p_s4_o23_0),
.I3(p_s4_o23_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER25////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo25 (
.O6(P[25]),
.O5(G[25]),
.I0(p_s4_o25_0),
.I1(p_s4_o25_1),
.I2(p_s4_o24_0),
.I3(p_s4_o24_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER26////////////

wire p_s4_o26_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o26_t264_z0_v0 (
.O6(p_s4_o26_1),
.O5(),
.I0(p_s3_o26_0),
.I1(p_s3_o26_1),
.I2(p_s3_o26_2),
.I3(p_s3_o26_3),
.I4(p_s2_o26_6),
.I5(p_s3_o27_0));

wire p_s4_o27_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o26_t264_z1_v0 (
.O6(p_s4_o27_0),
.O5(),
.I0(p_s3_o26_0),
.I1(p_s3_o26_1),
.I2(p_s3_o26_2),
.I3(p_s3_o26_3),
.I4(p_s2_o26_6),
.I5(p_s3_o27_0));

wire p_s4_o28_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o26_t264_z2_v0 (
.O6(p_s4_o28_0),
.O5(),
.I0(p_s3_o26_0),
.I1(p_s3_o26_1),
.I2(p_s3_o26_2),
.I3(p_s3_o26_3),
.I4(p_s2_o26_6),
.I5(p_s3_o27_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo26 (
.O6(P[26]),
.O5(G[26]),
.I0(p_s4_o26_0),
.I1(p_s4_o26_1),
.I2(p_s4_o25_0),
.I3(p_s4_o25_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER27////////////

wire p_s4_o28_1;
wire p_s4_o27_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o27_t276_z0_v0 (
.O6(p_s4_o28_1),
.O5(p_s4_o27_1),
.I0(p_s3_o27_1),
.I1(p_s3_o27_2),
.I2(p_s3_o27_3),
.I3(p_s3_o28_0),
.I4(p_s3_o28_1),
.I5(1'b1));

wire p_s4_o29_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o27_t276_z1_v0 (
.O6(p_s4_o29_0),
.O5(),
.I0(p_s3_o27_1),
.I1(p_s3_o27_2),
.I2(p_s3_o27_3),
.I3(p_s3_o28_0),
.I4(p_s3_o28_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo27 (
.O6(P[27]),
.O5(G[27]),
.I0(p_s4_o27_0),
.I1(p_s4_o27_1),
.I2(p_s4_o26_0),
.I3(p_s4_o26_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER28////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo28 (
.O6(P[28]),
.O5(G[28]),
.I0(p_s4_o28_0),
.I1(p_s4_o28_1),
.I2(p_s4_o27_0),
.I3(p_s4_o27_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER29////////////

wire p_s4_o30_0;
wire p_s4_o29_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o29_t277_z0_v0 (
.O6(p_s4_o30_0),
.O5(p_s4_o29_1),
.I0(p_s3_o29_0),
.I1(p_s3_o29_1),
.I2(p_s3_o29_2),
.I3(p_s3_o30_0),
.I4(p_s3_o30_1),
.I5(1'b1));

wire p_s4_o31_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o29_t277_z1_v0 (
.O6(p_s4_o31_0),
.O5(),
.I0(p_s3_o29_0),
.I1(p_s3_o29_1),
.I2(p_s3_o29_2),
.I3(p_s3_o30_0),
.I4(p_s3_o30_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo29 (
.O6(P[29]),
.O5(G[29]),
.I0(p_s4_o29_0),
.I1(p_s4_o29_1),
.I2(p_s4_o28_0),
.I3(p_s4_o28_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER30////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo30 (
.O6(P[30]),
.O5(G[30]),
.I0(p_s4_o30_0),
.I1(p_s3_o30_2),
.I2(p_s4_o29_0),
.I3(p_s4_o29_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER31////////////

wire p_s4_o32_0;
wire p_s4_o31_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o31_t278_z0_v0 (
.O6(p_s4_o32_0),
.O5(p_s4_o31_1),
.I0(p_s3_o31_0),
.I1(p_s3_o31_1),
.I2(p_s3_o31_2),
.I3(p_s3_o32_0),
.I4(p_s3_o32_1),
.I5(1'b1));

wire p_s4_o33_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o31_t278_z1_v0 (
.O6(p_s4_o33_0),
.O5(),
.I0(p_s3_o31_0),
.I1(p_s3_o31_1),
.I2(p_s3_o31_2),
.I3(p_s3_o32_0),
.I4(p_s3_o32_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo31 (
.O6(P[31]),
.O5(G[31]),
.I0(p_s4_o31_0),
.I1(p_s4_o31_1),
.I2(p_s4_o30_0),
.I3(p_s3_o30_2),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER32////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo32 (
.O6(P[32]),
.O5(G[32]),
.I0(p_s4_o32_0),
.I1(p_s3_o32_2),
.I2(p_s4_o31_0),
.I3(p_s4_o31_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER33////////////

wire p_s4_o33_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o33_t265_z0_v0 (
.O6(p_s4_o33_1),
.O5(),
.I0(p_s3_o33_0),
.I1(p_s3_o33_1),
.I2(p_s3_o33_2),
.I3(p_s2_o33_4),
.I4(p_s2_o33_5),
.I5(p_s3_o34_0));

wire p_s4_o34_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o33_t265_z1_v0 (
.O6(p_s4_o34_0),
.O5(),
.I0(p_s3_o33_0),
.I1(p_s3_o33_1),
.I2(p_s3_o33_2),
.I3(p_s2_o33_4),
.I4(p_s2_o33_5),
.I5(p_s3_o34_0));

wire p_s4_o35_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o33_t265_z2_v0 (
.O6(p_s4_o35_0),
.O5(),
.I0(p_s3_o33_0),
.I1(p_s3_o33_1),
.I2(p_s3_o33_2),
.I3(p_s2_o33_4),
.I4(p_s2_o33_5),
.I5(p_s3_o34_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo33 (
.O6(P[33]),
.O5(G[33]),
.I0(p_s4_o33_0),
.I1(p_s4_o33_1),
.I2(p_s4_o32_0),
.I3(p_s3_o32_2),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER34////////////

wire p_s4_o35_1;
wire p_s4_o34_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o34_t279_z0_v0 (
.O6(p_s4_o35_1),
.O5(p_s4_o34_1),
.I0(p_s3_o34_1),
.I1(p_s3_o34_2),
.I2(p_s2_o34_5),
.I3(p_s3_o35_0),
.I4(p_s3_o35_1),
.I5(1'b1));

wire p_s4_o36_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o34_t279_z1_v0 (
.O6(p_s4_o36_0),
.O5(),
.I0(p_s3_o34_1),
.I1(p_s3_o34_2),
.I2(p_s2_o34_5),
.I3(p_s3_o35_0),
.I4(p_s3_o35_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo34 (
.O6(P[34]),
.O5(G[34]),
.I0(p_s4_o34_0),
.I1(p_s4_o34_1),
.I2(p_s4_o33_0),
.I3(p_s4_o33_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER35////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo35 (
.O6(P[35]),
.O5(G[35]),
.I0(p_s4_o35_0),
.I1(p_s4_o35_1),
.I2(p_s4_o34_0),
.I3(p_s4_o34_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER36////////////

wire p_s4_o37_0;
wire p_s4_o36_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o36_t280_z0_v0 (
.O6(p_s4_o37_0),
.O5(p_s4_o36_1),
.I0(p_s3_o36_0),
.I1(p_s3_o36_1),
.I2(p_s3_o36_2),
.I3(p_s3_o37_0),
.I4(p_s3_o37_1),
.I5(1'b1));

wire p_s4_o38_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o36_t280_z1_v0 (
.O6(p_s4_o38_0),
.O5(),
.I0(p_s3_o36_0),
.I1(p_s3_o36_1),
.I2(p_s3_o36_2),
.I3(p_s3_o37_0),
.I4(p_s3_o37_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo36 (
.O6(P[36]),
.O5(G[36]),
.I0(p_s4_o36_0),
.I1(p_s4_o36_1),
.I2(p_s4_o35_0),
.I3(p_s4_o35_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER37////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo37 (
.O6(P[37]),
.O5(G[37]),
.I0(p_s4_o37_0),
.I1(p_s3_o37_2),
.I2(p_s4_o36_0),
.I3(p_s4_o36_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER38////////////

wire p_s4_o39_0;
wire p_s4_o38_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s4_o38_t251_z0_v0 (
.O6(p_s4_o39_0),
.O5(p_s4_o38_1),
.I0(p_s3_o38_0),
.I1(p_s3_o38_1),
.I2(p_s3_o38_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo38 (
.O6(P[38]),
.O5(G[38]),
.I0(p_s4_o38_0),
.I1(p_s4_o38_1),
.I2(p_s4_o37_0),
.I3(p_s3_o37_2),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER39////////////

wire p_s4_o39_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o39_t266_z0_v0 (
.O6(p_s4_o39_1),
.O5(),
.I0(p_s3_o39_0),
.I1(p_s3_o39_1),
.I2(p_s3_o39_2),
.I3(p_s2_o39_4),
.I4(p_s2_o39_5),
.I5(p_s3_o40_0));

wire p_s4_o40_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o39_t266_z1_v0 (
.O6(p_s4_o40_0),
.O5(),
.I0(p_s3_o39_0),
.I1(p_s3_o39_1),
.I2(p_s3_o39_2),
.I3(p_s2_o39_4),
.I4(p_s2_o39_5),
.I5(p_s3_o40_0));

wire p_s4_o41_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o39_t266_z2_v0 (
.O6(p_s4_o41_0),
.O5(),
.I0(p_s3_o39_0),
.I1(p_s3_o39_1),
.I2(p_s3_o39_2),
.I3(p_s2_o39_4),
.I4(p_s2_o39_5),
.I5(p_s3_o40_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo39 (
.O6(P[39]),
.O5(G[39]),
.I0(p_s4_o39_0),
.I1(p_s4_o39_1),
.I2(p_s4_o38_0),
.I3(p_s4_o38_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER40////////////

wire p_s4_o41_1;
wire p_s4_o40_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o40_t281_z0_v0 (
.O6(p_s4_o41_1),
.O5(p_s4_o40_1),
.I0(p_s3_o40_1),
.I1(p_s3_o40_2),
.I2(p_s2_o40_5),
.I3(p_s3_o41_0),
.I4(p_s3_o41_1),
.I5(1'b1));

wire p_s4_o42_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o40_t281_z1_v0 (
.O6(p_s4_o42_0),
.O5(),
.I0(p_s3_o40_1),
.I1(p_s3_o40_2),
.I2(p_s2_o40_5),
.I3(p_s3_o41_0),
.I4(p_s3_o41_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo40 (
.O6(P[40]),
.O5(G[40]),
.I0(p_s4_o40_0),
.I1(p_s4_o40_1),
.I2(p_s4_o39_0),
.I3(p_s4_o39_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER41////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo41 (
.O6(P[41]),
.O5(G[41]),
.I0(p_s4_o41_0),
.I1(p_s4_o41_1),
.I2(p_s4_o40_0),
.I3(p_s4_o40_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER42////////////

wire p_s4_o42_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o42_t267_z0_v0 (
.O6(p_s4_o42_1),
.O5(),
.I0(p_s3_o42_0),
.I1(p_s3_o42_1),
.I2(p_s3_o42_2),
.I3(p_s2_o42_4),
.I4(p_s2_o42_5),
.I5(p_s3_o43_0));

wire p_s4_o43_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o42_t267_z1_v0 (
.O6(p_s4_o43_0),
.O5(),
.I0(p_s3_o42_0),
.I1(p_s3_o42_1),
.I2(p_s3_o42_2),
.I3(p_s2_o42_4),
.I4(p_s2_o42_5),
.I5(p_s3_o43_0));

wire p_s4_o44_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o42_t267_z2_v0 (
.O6(p_s4_o44_0),
.O5(),
.I0(p_s3_o42_0),
.I1(p_s3_o42_1),
.I2(p_s3_o42_2),
.I3(p_s2_o42_4),
.I4(p_s2_o42_5),
.I5(p_s3_o43_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo42 (
.O6(P[42]),
.O5(G[42]),
.I0(p_s4_o42_0),
.I1(p_s4_o42_1),
.I2(p_s4_o41_0),
.I3(p_s4_o41_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER43////////////

wire p_s4_o44_1;
wire p_s4_o43_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o43_t282_z0_v0 (
.O6(p_s4_o44_1),
.O5(p_s4_o43_1),
.I0(p_s3_o43_1),
.I1(p_s3_o43_2),
.I2(p_s2_o43_5),
.I3(p_s3_o44_0),
.I4(p_s3_o44_1),
.I5(1'b1));

wire p_s4_o45_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o43_t282_z1_v0 (
.O6(p_s4_o45_0),
.O5(),
.I0(p_s3_o43_1),
.I1(p_s3_o43_2),
.I2(p_s2_o43_5),
.I3(p_s3_o44_0),
.I4(p_s3_o44_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo43 (
.O6(P[43]),
.O5(G[43]),
.I0(p_s4_o43_0),
.I1(p_s4_o43_1),
.I2(p_s4_o42_0),
.I3(p_s4_o42_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER44////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo44 (
.O6(P[44]),
.O5(G[44]),
.I0(p_s4_o44_0),
.I1(p_s4_o44_1),
.I2(p_s4_o43_0),
.I3(p_s4_o43_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER45////////////

wire p_s4_o46_0;
wire p_s4_o45_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o45_t283_z0_v0 (
.O6(p_s4_o46_0),
.O5(p_s4_o45_1),
.I0(p_s3_o45_0),
.I1(p_s3_o45_1),
.I2(p_s3_o45_2),
.I3(p_s3_o46_0),
.I4(p_s3_o46_1),
.I5(1'b1));

wire p_s4_o47_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o45_t283_z1_v0 (
.O6(p_s4_o47_0),
.O5(),
.I0(p_s3_o45_0),
.I1(p_s3_o45_1),
.I2(p_s3_o45_2),
.I3(p_s3_o46_0),
.I4(p_s3_o46_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo45 (
.O6(P[45]),
.O5(G[45]),
.I0(p_s4_o45_0),
.I1(p_s4_o45_1),
.I2(p_s4_o44_0),
.I3(p_s4_o44_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER46////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo46 (
.O6(P[46]),
.O5(G[46]),
.I0(p_s4_o46_0),
.I1(p_s3_o46_2),
.I2(p_s4_o45_0),
.I3(p_s4_o45_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER47////////////

wire p_s4_o47_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o47_t268_z0_v0 (
.O6(p_s4_o47_1),
.O5(),
.I0(p_s3_o47_0),
.I1(p_s3_o47_1),
.I2(p_s3_o47_2),
.I3(p_s3_o47_3),
.I4(p_s1_o47_5),
.I5(p_s3_o48_0));

wire p_s4_o48_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o47_t268_z1_v0 (
.O6(p_s4_o48_0),
.O5(),
.I0(p_s3_o47_0),
.I1(p_s3_o47_1),
.I2(p_s3_o47_2),
.I3(p_s3_o47_3),
.I4(p_s1_o47_5),
.I5(p_s3_o48_0));

wire p_s4_o49_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o47_t268_z2_v0 (
.O6(p_s4_o49_0),
.O5(),
.I0(p_s3_o47_0),
.I1(p_s3_o47_1),
.I2(p_s3_o47_2),
.I3(p_s3_o47_3),
.I4(p_s1_o47_5),
.I5(p_s3_o48_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo47 (
.O6(P[47]),
.O5(G[47]),
.I0(p_s4_o47_0),
.I1(p_s4_o47_1),
.I2(p_s4_o46_0),
.I3(p_s3_o46_2),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER48////////////

wire p_s4_o49_1;
wire p_s4_o48_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o48_t284_z0_v0 (
.O6(p_s4_o49_1),
.O5(p_s4_o48_1),
.I0(p_s3_o48_1),
.I1(p_s3_o48_2),
.I2(p_s3_o48_3),
.I3(p_s3_o49_0),
.I4(p_s3_o49_1),
.I5(1'b1));

wire p_s4_o50_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o48_t284_z1_v0 (
.O6(p_s4_o50_0),
.O5(),
.I0(p_s3_o48_1),
.I1(p_s3_o48_2),
.I2(p_s3_o48_3),
.I3(p_s3_o49_0),
.I4(p_s3_o49_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo48 (
.O6(P[48]),
.O5(G[48]),
.I0(p_s4_o48_0),
.I1(p_s4_o48_1),
.I2(p_s4_o47_0),
.I3(p_s4_o47_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER49////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo49 (
.O6(P[49]),
.O5(G[49]),
.I0(p_s4_o49_0),
.I1(p_s4_o49_1),
.I2(p_s4_o48_0),
.I3(p_s4_o48_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER50////////////

wire p_s4_o50_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o50_t269_z0_v0 (
.O6(p_s4_o50_1),
.O5(),
.I0(p_s3_o50_0),
.I1(p_s3_o50_1),
.I2(p_s3_o50_2),
.I3(p_s3_o50_3),
.I4(p_s2_o50_6),
.I5(p_s3_o51_0));

wire p_s4_o51_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o50_t269_z1_v0 (
.O6(p_s4_o51_0),
.O5(),
.I0(p_s3_o50_0),
.I1(p_s3_o50_1),
.I2(p_s3_o50_2),
.I3(p_s3_o50_3),
.I4(p_s2_o50_6),
.I5(p_s3_o51_0));

wire p_s4_o52_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o50_t269_z2_v0 (
.O6(p_s4_o52_0),
.O5(),
.I0(p_s3_o50_0),
.I1(p_s3_o50_1),
.I2(p_s3_o50_2),
.I3(p_s3_o50_3),
.I4(p_s2_o50_6),
.I5(p_s3_o51_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo50 (
.O6(P[50]),
.O5(G[50]),
.I0(p_s4_o50_0),
.I1(p_s4_o50_1),
.I2(p_s4_o49_0),
.I3(p_s4_o49_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER51////////////

wire p_s4_o52_1;
wire p_s4_o51_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o51_t285_z0_v0 (
.O6(p_s4_o52_1),
.O5(p_s4_o51_1),
.I0(p_s3_o51_1),
.I1(p_s3_o51_2),
.I2(p_s3_o51_3),
.I3(p_s3_o52_0),
.I4(p_s3_o52_1),
.I5(1'b1));

wire p_s4_o53_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o51_t285_z1_v0 (
.O6(p_s4_o53_0),
.O5(),
.I0(p_s3_o51_1),
.I1(p_s3_o51_2),
.I2(p_s3_o51_3),
.I3(p_s3_o52_0),
.I4(p_s3_o52_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo51 (
.O6(P[51]),
.O5(G[51]),
.I0(p_s4_o51_0),
.I1(p_s4_o51_1),
.I2(p_s4_o50_0),
.I3(p_s4_o50_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER52////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo52 (
.O6(P[52]),
.O5(G[52]),
.I0(p_s4_o52_0),
.I1(p_s4_o52_1),
.I2(p_s4_o51_0),
.I3(p_s4_o51_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER53////////////

wire p_s4_o53_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o53_t270_z0_v0 (
.O6(p_s4_o53_1),
.O5(),
.I0(p_s3_o53_0),
.I1(p_s3_o53_1),
.I2(p_s3_o53_2),
.I3(p_s3_o53_3),
.I4(p_s3_o53_4),
.I5(p_s3_o54_0));

wire p_s4_o54_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o53_t270_z1_v0 (
.O6(p_s4_o54_0),
.O5(),
.I0(p_s3_o53_0),
.I1(p_s3_o53_1),
.I2(p_s3_o53_2),
.I3(p_s3_o53_3),
.I4(p_s3_o53_4),
.I5(p_s3_o54_0));

wire p_s4_o55_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o53_t270_z2_v0 (
.O6(p_s4_o55_0),
.O5(),
.I0(p_s3_o53_0),
.I1(p_s3_o53_1),
.I2(p_s3_o53_2),
.I3(p_s3_o53_3),
.I4(p_s3_o53_4),
.I5(p_s3_o54_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo53 (
.O6(P[53]),
.O5(G[53]),
.I0(p_s4_o53_0),
.I1(p_s4_o53_1),
.I2(p_s4_o52_0),
.I3(p_s4_o52_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER54////////////

wire p_s4_o55_1;
wire p_s4_o54_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o54_t286_z0_v0 (
.O6(p_s4_o55_1),
.O5(p_s4_o54_1),
.I0(p_s3_o54_1),
.I1(p_s3_o54_2),
.I2(p_s3_o54_3),
.I3(p_s3_o55_0),
.I4(p_s3_o55_1),
.I5(1'b1));

wire p_s4_o56_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o54_t286_z1_v0 (
.O6(p_s4_o56_0),
.O5(),
.I0(p_s3_o54_1),
.I1(p_s3_o54_2),
.I2(p_s3_o54_3),
.I3(p_s3_o55_0),
.I4(p_s3_o55_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo54 (
.O6(P[54]),
.O5(G[54]),
.I0(p_s4_o54_0),
.I1(p_s4_o54_1),
.I2(p_s4_o53_0),
.I3(p_s4_o53_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER55////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo55 (
.O6(P[55]),
.O5(G[55]),
.I0(p_s4_o55_0),
.I1(p_s4_o55_1),
.I2(p_s4_o54_0),
.I3(p_s4_o54_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER56////////////

wire p_s4_o57_0;
wire p_s4_o56_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s4_o56_t252_z0_v0 (
.O6(p_s4_o57_0),
.O5(p_s4_o56_1),
.I0(p_s3_o56_0),
.I1(p_s3_o56_1),
.I2(p_s2_o56_1),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo56 (
.O6(P[56]),
.O5(G[56]),
.I0(p_s4_o56_0),
.I1(p_s4_o56_1),
.I2(p_s4_o55_0),
.I3(p_s4_o55_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER57////////////

wire p_s4_o58_0;
wire p_s4_o57_1;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s4_o57_t253_z0_v0 (
.O6(p_s4_o58_0),
.O5(p_s4_o57_1),
.I0(a[29]),
.I1(b[31]),
.I2(p_s3_o57_0),
.I3(p_s3_o57_1),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo57 (
.O6(P[57]),
.O5(G[57]),
.I0(p_s4_o57_0),
.I1(p_s4_o57_1),
.I2(p_s4_o56_0),
.I3(p_s4_o56_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER58////////////

wire p_s4_o59_0;
wire p_s4_o58_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s4_o58_t254_z0_v0 (
.O6(p_s4_o59_0),
.O5(p_s4_o58_1),
.I0(a[31]),
.I1(b[30]),
.I2(a[30]),
.I3(b[31]),
.I4(p_s3_o58_0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo58 (
.O6(P[58]),
.O5(G[58]),
.I0(p_s4_o58_0),
.I1(p_s4_o58_1),
.I2(p_s4_o57_0),
.I3(p_s4_o57_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER59////////////

LUT6_2 #(
.INIT(64'h87777888F8888000)
) LUT6_2_inst_ooo (
.O6(P[59]),
.O5(G[59]),
.I0(b[31]),
.I1(a[31]),
.I2(p_s4_o58_0),
.I3(p_s4_o58_1),
.I4(p_s4_o59_0),
.I5(1'b1));

wire [3:0] carry_o_0;
CARRY4  CARRY4_inst_0(
.CO(carry_o_0),
.O(r[6:3]),
.CI(C1),
.CYINIT(1'b0),
.DI(G[3:0]),
.S(P[3:0]));

wire [3:0] carry_o_1;
CARRY4  CARRY4_inst_1(
.CO(carry_o_1),
.O(r[10:7]),
.CI(carry_o_0[3]),
.CYINIT(1'b0),
.DI(G[7:4]),
.S(P[7:4]));

wire [3:0] carry_o_2;
CARRY4  CARRY4_inst_2(
.CO(carry_o_2),
.O(r[14:11]),
.CI(carry_o_1[3]),
.CYINIT(1'b0),
.DI(G[11:8]),
.S(P[11:8]));

wire [3:0] carry_o_3;
CARRY4  CARRY4_inst_3(
.CO(carry_o_3),
.O(r[18:15]),
.CI(carry_o_2[3]),
.CYINIT(1'b0),
.DI(G[15:12]),
.S(P[15:12]));

wire [3:0] carry_o_4;
CARRY4  CARRY4_inst_4(
.CO(carry_o_4),
.O(r[22:19]),
.CI(carry_o_3[3]),
.CYINIT(1'b0),
.DI(G[19:16]),
.S(P[19:16]));

wire [3:0] carry_o_5;
CARRY4  CARRY4_inst_5(
.CO(carry_o_5),
.O(r[26:23]),
.CI(carry_o_4[3]),
.CYINIT(1'b0),
.DI(G[23:20]),
.S(P[23:20]));

wire [3:0] carry_o_6;
CARRY4  CARRY4_inst_6(
.CO(carry_o_6),
.O(r[30:27]),
.CI(carry_o_5[3]),
.CYINIT(1'b0),
.DI(G[27:24]),
.S(P[27:24]));

wire [3:0] carry_o_7;
CARRY4  CARRY4_inst_7(
.CO(carry_o_7),
.O(r[34:31]),
.CI(carry_o_6[3]),
.CYINIT(1'b0),
.DI(G[31:28]),
.S(P[31:28]));

wire [3:0] carry_o_8;
CARRY4  CARRY4_inst_8(
.CO(carry_o_8),
.O(r[38:35]),
.CI(carry_o_7[3]),
.CYINIT(1'b0),
.DI(G[35:32]),
.S(P[35:32]));

wire [3:0] carry_o_9;
CARRY4  CARRY4_inst_9(
.CO(carry_o_9),
.O(r[42:39]),
.CI(carry_o_8[3]),
.CYINIT(1'b0),
.DI(G[39:36]),
.S(P[39:36]));

wire [3:0] carry_o_10;
CARRY4  CARRY4_inst_10(
.CO(carry_o_10),
.O(r[46:43]),
.CI(carry_o_9[3]),
.CYINIT(1'b0),
.DI(G[43:40]),
.S(P[43:40]));

wire [3:0] carry_o_11;
CARRY4  CARRY4_inst_11(
.CO(carry_o_11),
.O(r[50:47]),
.CI(carry_o_10[3]),
.CYINIT(1'b0),
.DI(G[47:44]),
.S(P[47:44]));

wire [3:0] carry_o_12;
CARRY4  CARRY4_inst_12(
.CO(carry_o_12),
.O(r[54:51]),
.CI(carry_o_11[3]),
.CYINIT(1'b0),
.DI(G[51:48]),
.S(P[51:48]));

wire [3:0] carry_o_13;
CARRY4  CARRY4_inst_13(
.CO(carry_o_13),
.O(r[58:55]),
.CI(carry_o_12[3]),
.CYINIT(1'b0),
.DI(G[55:52]),
.S(P[55:52]));

wire [3:0] carry_o_14;
CARRY4  CARRY4_inst_14(
.CO(carry_o_14),
.O(r[62:59]),
.CI(carry_o_13[3]),
.CYINIT(1'b0),
.DI(G[59:56]),
.S(P[59:56]));

assign  r[63] = carry_o_14[3] | (P[59] & G[59]);
//v2024-09-17 10:16:39.991458
endmodule

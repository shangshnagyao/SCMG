module mult_8b_5s ( 
input [8-1:0] a,
input [8-1:0] b,
output [2*8-1:0] r
);

// Target value:54
wire [11:0] P;
wire [11:0] G;

// 4 normal LUT
LUT6_2 #(
.INIT(64'h78887888C0C0C0C0)
) LUT6_2_inst_f0 (
.O6(r[1]),
.O5(r[0]),
.I0(b[1]),
.I1(a[0]),
.I2(b[0]),
.I3(a[1]),
.I4(1'b1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h47777888B8887888)
) LUT6_2_inst_f1 (
.O6(r[2]),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

LUT6_2 #(
.INIT(64'hF8888000C0008000)
) LUT6_2_inst_f2 (
.O6(C1),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

LUT6_2 #(
.INIT(64'h8000000000000000)
) LUT6_2_inst_f3 (
.O6(C0),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

/////////STEP0----ORDER0////////////

wire p_s0_o0_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o0_t0_z0_v0 (
.O6(p_s0_o0_0),
.O5(),
.I0(a[3]),
.I1(b[0]),
.I2(a[2]),
.I3(b[1]),
.I4(a[1]),
.I5(b[2]));

wire p_s0_o1_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o0_t0_z1_v0 (
.O6(p_s0_o1_0),
.O5(),
.I0(a[3]),
.I1(b[0]),
.I2(a[2]),
.I3(b[1]),
.I4(a[1]),
.I5(b[2]));

/////////STEP0----ORDER1////////////

/////////STEP0----ORDER2////////////

/////////STEP0----ORDER3////////////

wire p_s0_o3_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o3_t1_z0_v0 (
.O6(p_s0_o3_0),
.O5(),
.I0(a[6]),
.I1(b[0]),
.I2(a[5]),
.I3(b[1]),
.I4(a[4]),
.I5(b[2]));

wire p_s0_o4_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o3_t1_z1_v0 (
.O6(p_s0_o4_0),
.O5(),
.I0(a[6]),
.I1(b[0]),
.I2(a[5]),
.I3(b[1]),
.I4(a[4]),
.I5(b[2]));

/////////STEP0----ORDER4////////////

/////////STEP0----ORDER5////////////

/////////STEP0----ORDER6////////////

wire p_s0_o6_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o6_t2_z0_v0 (
.O6(p_s0_o6_0),
.O5(),
.I0(a[7]),
.I1(b[2]),
.I2(a[6]),
.I3(b[3]),
.I4(a[5]),
.I5(b[4]));

wire p_s0_o7_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o6_t2_z1_v0 (
.O6(p_s0_o7_0),
.O5(),
.I0(a[7]),
.I1(b[2]),
.I2(a[6]),
.I3(b[3]),
.I4(a[5]),
.I5(b[4]));

/////////STEP0----ORDER7////////////

/////////STEP0----ORDER8////////////

/////////STEP0----ORDER9////////////

/////////STEP0----ORDER10////////////

/////////STEP0----ORDER11////////////

/////////STEP1----ORDER0////////////

/////////STEP1----ORDER1////////////

wire p_s1_o2_0;
wire p_s1_o1_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o1_t3_z0_v0 (
.O6(p_s1_o2_0),
.O5(p_s1_o1_0),
.I0(a[4]),
.I1(b[0]),
.I2(a[3]),
.I3(b[1]),
.I4(p_s0_o1_0),
.I5(1'b1));

/////////STEP1----ORDER2////////////

/////////STEP1----ORDER3////////////

wire p_s1_o4_0;
wire p_s1_o3_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o3_t4_z0_v0 (
.O6(p_s1_o4_0),
.O5(p_s1_o3_0),
.I0(a[3]),
.I1(b[3]),
.I2(a[2]),
.I3(b[4]),
.I4(p_s0_o3_0),
.I5(1'b1));

/////////STEP1----ORDER4////////////

wire p_s1_o5_0;
wire p_s1_o4_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o4_t5_z0_v0 (
.O6(p_s1_o5_0),
.O5(p_s1_o4_1),
.I0(a[7]),
.I1(b[0]),
.I2(a[6]),
.I3(b[1]),
.I4(p_s0_o4_0),
.I5(1'b1));

/////////STEP1----ORDER5////////////

/////////STEP1----ORDER6////////////

/////////STEP1----ORDER7////////////

wire p_s1_o8_0;
wire p_s1_o7_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o7_t6_z0_v0 (
.O6(p_s1_o8_0),
.O5(p_s1_o7_0),
.I0(a[7]),
.I1(b[3]),
.I2(a[6]),
.I3(b[4]),
.I4(p_s0_o7_0),
.I5(1'b1));

/////////STEP1----ORDER8////////////

/////////STEP1----ORDER9////////////

/////////STEP1----ORDER10////////////

/////////STEP1----ORDER11////////////

/////////STEP2----ORDER0////////////

/////////STEP2----ORDER1////////////

wire p_s2_o2_0;
wire p_s2_o1_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o1_t7_z0_v0 (
.O6(p_s2_o2_0),
.O5(p_s2_o1_0),
.I0(a[2]),
.I1(b[2]),
.I2(a[1]),
.I3(b[3]),
.I4(p_s1_o1_0),
.I5(1'b1));

/////////STEP2----ORDER2////////////

wire p_s2_o3_0;
wire p_s2_o2_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o2_t8_z0_v0 (
.O6(p_s2_o3_0),
.O5(p_s2_o2_1),
.I0(a[5]),
.I1(b[0]),
.I2(a[4]),
.I3(b[1]),
.I4(p_s1_o2_0),
.I5(1'b1));

/////////STEP2----ORDER3////////////

wire p_s2_o4_0;
wire p_s2_o3_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o3_t9_z0_v0 (
.O6(p_s2_o4_0),
.O5(p_s2_o3_1),
.I0(a[1]),
.I1(b[5]),
.I2(a[0]),
.I3(b[6]),
.I4(p_s1_o3_0),
.I5(1'b1));

/////////STEP2----ORDER4////////////

wire p_s2_o5_0;
wire p_s2_o4_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o4_t10_z0_v0 (
.O6(p_s2_o5_0),
.O5(p_s2_o4_1),
.I0(a[5]),
.I1(b[2]),
.I2(a[4]),
.I3(b[3]),
.I4(p_s1_o4_0),
.I5(1'b1));

wire p_s2_o5_1;
wire p_s2_o4_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o4_t10_z0_v1 (
.O6(p_s2_o5_1),
.O5(p_s2_o4_2),
.I0(a[3]),
.I1(b[4]),
.I2(a[2]),
.I3(b[5]),
.I4(p_s1_o4_1),
.I5(1'b1));

/////////STEP2----ORDER5////////////

wire p_s2_o6_0;
wire p_s2_o5_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o5_t11_z0_v0 (
.O6(p_s2_o6_0),
.O5(p_s2_o5_2),
.I0(a[7]),
.I1(b[1]),
.I2(a[6]),
.I3(b[2]),
.I4(p_s1_o5_0),
.I5(1'b1));

/////////STEP2----ORDER6////////////

wire p_s2_o7_0;
wire p_s2_o6_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o6_t12_z0_v0 (
.O6(p_s2_o7_0),
.O5(p_s2_o6_1),
.I0(a[4]),
.I1(b[5]),
.I2(a[3]),
.I3(b[6]),
.I4(p_s0_o6_0),
.I5(1'b1));

/////////STEP2----ORDER7////////////

wire p_s2_o8_0;
wire p_s2_o7_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o7_t13_z0_v0 (
.O6(p_s2_o8_0),
.O5(p_s2_o7_1),
.I0(a[5]),
.I1(b[5]),
.I2(a[4]),
.I3(b[6]),
.I4(p_s1_o7_0),
.I5(1'b1));

/////////STEP2----ORDER8////////////

wire p_s2_o9_0;
wire p_s2_o8_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o8_t14_z0_v0 (
.O6(p_s2_o9_0),
.O5(p_s2_o8_1),
.I0(a[7]),
.I1(b[4]),
.I2(a[6]),
.I3(b[5]),
.I4(p_s1_o8_0),
.I5(1'b1));

/////////STEP2----ORDER9////////////

/////////STEP2----ORDER10////////////

/////////STEP2----ORDER11////////////

/////////STEP3----ORDER0////////////

/////////STEP3----ORDER1////////////

/////////STEP3----ORDER2////////////

wire p_s3_o3_0;
wire p_s3_o2_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o2_t18_z0_v0 (
.O6(p_s3_o3_0),
.O5(p_s3_o2_0),
.I0(a[3]),
.I1(b[2]),
.I2(a[2]),
.I3(b[3]),
.I4(p_s2_o2_0),
.I5(1'b1));

wire p_s3_o3_1;
wire p_s3_o2_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o2_t18_z0_v1 (
.O6(p_s3_o3_1),
.O5(p_s3_o2_1),
.I0(a[1]),
.I1(b[4]),
.I2(a[0]),
.I3(b[5]),
.I4(p_s2_o2_1),
.I5(1'b1));

/////////STEP3----ORDER3////////////

/////////STEP3----ORDER4////////////

wire p_s3_o5_0;
wire p_s3_o4_0;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o4_t15_z0_v0 (
.O6(p_s3_o5_0),
.O5(p_s3_o4_0),
.I0(p_s2_o4_0),
.I1(p_s2_o4_1),
.I2(p_s2_o4_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER5////////////

wire p_s3_o6_0;
wire p_s3_o5_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o5_t19_z0_v0 (
.O6(p_s3_o6_0),
.O5(p_s3_o5_1),
.I0(a[5]),
.I1(b[3]),
.I2(a[4]),
.I3(b[4]),
.I4(p_s2_o5_0),
.I5(1'b1));

wire p_s3_o6_1;
wire p_s3_o5_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o5_t19_z0_v1 (
.O6(p_s3_o6_1),
.O5(p_s3_o5_2),
.I0(a[3]),
.I1(b[5]),
.I2(a[2]),
.I3(b[6]),
.I4(p_s2_o5_1),
.I5(1'b1));

wire p_s3_o6_2;
wire p_s3_o5_3;
LUT6_2 #(
.INIT(64'h8080808078787878)
) LUT6_2_inst_s3_o5_t22_z0_v0 (
.O6(p_s3_o6_2),
.O5(p_s3_o5_3),
.I0(a[1]),
.I1(b[7]),
.I2(p_s2_o5_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER6////////////

wire p_s3_o7_0;
wire p_s3_o6_3;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o6_t16_z0_v0 (
.O6(p_s3_o7_0),
.O5(p_s3_o6_3),
.I0(a[2]),
.I1(b[7]),
.I2(p_s2_o6_0),
.I3(p_s2_o6_1),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER7////////////

wire p_s3_o8_0;
wire p_s3_o7_1;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o7_t17_z0_v0 (
.O6(p_s3_o8_0),
.O5(p_s3_o7_1),
.I0(a[3]),
.I1(b[7]),
.I2(p_s2_o7_0),
.I3(p_s2_o7_1),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER8////////////

wire p_s3_o9_0;
wire p_s3_o8_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o8_t20_z0_v0 (
.O6(p_s3_o9_0),
.O5(p_s3_o8_1),
.I0(a[5]),
.I1(b[6]),
.I2(a[4]),
.I3(b[7]),
.I4(p_s2_o8_0),
.I5(1'b1));

/////////STEP3----ORDER9////////////

wire p_s3_o10_0;
wire p_s3_o9_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o9_t21_z0_v0 (
.O6(p_s3_o10_0),
.O5(p_s3_o9_1),
.I0(a[7]),
.I1(b[5]),
.I2(a[6]),
.I3(b[6]),
.I4(p_s2_o9_0),
.I5(1'b1));

/////////STEP3----ORDER10////////////

/////////STEP3----ORDER11////////////

/////////STEP4----ORDER0////////////

LUT6_2 #(
.INIT(64'h8778877808800880)
) LUT6_2_inst_oo0 (
.O6(P[0]),
.O5(G[0]),
.I0(a[0]),
.I1(b[3]),
.I2(C0),
.I3(p_s0_o0_0),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER1////////////

LUT6_2 #(
.INIT(64'h8778787878000000)
) LUT6_2_inst_oo1 (
.O6(P[1]),
.O5(G[1]),
.I0(a[0]),
.I1(b[4]),
.I2(p_s2_o1_0),
.I3(C0),
.I4(p_s0_o0_0),
.I5(1'b1));

/////////STEP4----ORDER2////////////

LUT6_2 #(
.INIT(64'h9666666660000000)
) LUT6_2_inst_oo2 (
.O6(P[2]),
.O5(G[2]),
.I0(p_s3_o2_0),
.I1(p_s3_o2_1),
.I2(a[0]),
.I3(b[4]),
.I4(p_s2_o1_0),
.I5(1'b1));

/////////STEP4----ORDER3////////////

wire p_s4_o4_0;
wire p_s4_o3_0;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s4_o3_t23_z0_v0 (
.O6(p_s4_o4_0),
.O5(p_s4_o3_0),
.I0(p_s3_o3_0),
.I1(p_s3_o3_1),
.I2(p_s2_o3_0),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo3 (
.O6(P[3]),
.O5(G[3]),
.I0(p_s4_o3_0),
.I1(p_s2_o3_1),
.I2(p_s3_o2_0),
.I3(p_s3_o2_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER4////////////

wire p_s4_o5_0;
wire p_s4_o4_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s4_o4_t26_z0_v0 (
.O6(p_s4_o5_0),
.O5(p_s4_o4_1),
.I0(a[1]),
.I1(b[6]),
.I2(a[0]),
.I3(b[7]),
.I4(p_s3_o4_0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo4 (
.O6(P[4]),
.O5(G[4]),
.I0(p_s4_o4_0),
.I1(p_s4_o4_1),
.I2(p_s4_o3_0),
.I3(p_s2_o3_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER5////////////

wire p_s4_o6_0;
wire p_s4_o5_1;
LUT6_2 #(
.INIT(64'h81177EE869966996)
) LUT6_2_inst_s4_o5_t28_z0_v0 (
.O6(p_s4_o6_0),
.O5(p_s4_o5_1),
.I0(p_s3_o5_0),
.I1(p_s3_o5_1),
.I2(p_s3_o5_2),
.I3(p_s3_o5_3),
.I4(p_s3_o6_0),
.I5(1'b1));

wire p_s4_o7_0;
LUT6_2 #(
.INIT(64'hFEE88000FEE88000)
) LUT6_2_inst_s4_o5_t28_z1_v0 (
.O6(p_s4_o7_0),
.O5(),
.I0(p_s3_o5_0),
.I1(p_s3_o5_1),
.I2(p_s3_o5_2),
.I3(p_s3_o5_3),
.I4(p_s3_o6_0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo5 (
.O6(P[5]),
.O5(G[5]),
.I0(p_s4_o5_0),
.I1(p_s4_o5_1),
.I2(p_s4_o4_0),
.I3(p_s4_o4_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER6////////////

wire p_s4_o7_1;
wire p_s4_o6_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o6_t29_z0_v0 (
.O6(p_s4_o7_1),
.O5(p_s4_o6_1),
.I0(p_s3_o6_1),
.I1(p_s3_o6_2),
.I2(p_s3_o6_3),
.I3(p_s3_o7_0),
.I4(p_s3_o7_1),
.I5(1'b1));

wire p_s4_o8_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o6_t29_z1_v0 (
.O6(p_s4_o8_0),
.O5(),
.I0(p_s3_o6_1),
.I1(p_s3_o6_2),
.I2(p_s3_o6_3),
.I3(p_s3_o7_0),
.I4(p_s3_o7_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo6 (
.O6(P[6]),
.O5(G[6]),
.I0(p_s4_o6_0),
.I1(p_s4_o6_1),
.I2(p_s4_o5_0),
.I3(p_s4_o5_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER7////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo7 (
.O6(P[7]),
.O5(G[7]),
.I0(p_s4_o7_0),
.I1(p_s4_o7_1),
.I2(p_s4_o6_0),
.I3(p_s4_o6_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER8////////////

wire p_s4_o9_0;
wire p_s4_o8_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s4_o8_t24_z0_v0 (
.O6(p_s4_o9_0),
.O5(p_s4_o8_1),
.I0(p_s3_o8_0),
.I1(p_s3_o8_1),
.I2(p_s2_o8_1),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo8 (
.O6(P[8]),
.O5(G[8]),
.I0(p_s4_o8_0),
.I1(p_s4_o8_1),
.I2(p_s4_o7_0),
.I3(p_s4_o7_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER9////////////

wire p_s4_o10_0;
wire p_s4_o9_1;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s4_o9_t25_z0_v0 (
.O6(p_s4_o10_0),
.O5(p_s4_o9_1),
.I0(a[5]),
.I1(b[7]),
.I2(p_s3_o9_0),
.I3(p_s3_o9_1),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo9 (
.O6(P[9]),
.O5(G[9]),
.I0(p_s4_o9_0),
.I1(p_s4_o9_1),
.I2(p_s4_o8_0),
.I3(p_s4_o8_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER10////////////

wire p_s4_o11_0;
wire p_s4_o10_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s4_o10_t27_z0_v0 (
.O6(p_s4_o11_0),
.O5(p_s4_o10_1),
.I0(a[7]),
.I1(b[6]),
.I2(a[6]),
.I3(b[7]),
.I4(p_s3_o10_0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo10 (
.O6(P[10]),
.O5(G[10]),
.I0(p_s4_o10_0),
.I1(p_s4_o10_1),
.I2(p_s4_o9_0),
.I3(p_s4_o9_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER11////////////

LUT6_2 #(
.INIT(64'h87777888F8888000)
) LUT6_2_inst_ooo (
.O6(P[11]),
.O5(G[11]),
.I0(b[7]),
.I1(a[7]),
.I2(p_s4_o10_0),
.I3(p_s4_o10_1),
.I4(p_s4_o11_0),
.I5(1'b1));

wire [3:0] carry_o_0;
CARRY4  CARRY4_inst_0(
.CO(carry_o_0),
.O(r[6:3]),
.CI(C1),
.CYINIT(1'b0),
.DI(G[3:0]),
.S(P[3:0]));

wire [3:0] carry_o_1;
CARRY4  CARRY4_inst_1(
.CO(carry_o_1),
.O(r[10:7]),
.CI(carry_o_0[3]),
.CYINIT(1'b0),
.DI(G[7:4]),
.S(P[7:4]));

wire [3:0] carry_o_2;
CARRY4  CARRY4_inst_2(
.CO(carry_o_2),
.O(r[14:11]),
.CI(carry_o_1[3]),
.CYINIT(1'b0),
.DI(G[11:8]),
.S(P[11:8]));

assign  r[15] = carry_o_2[3] | (P[11] & G[11]);
//v2024-10-07 20:38:51.347707
endmodule

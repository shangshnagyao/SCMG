module mult_16b_5s ( 
input [16-1:0] a,
input [16-1:0] b,
output [2*16-1:0] r
);

// Target value:247
wire [27:0] P;
wire [27:0] G;

// 4 normal LUT
LUT6_2 #(
.INIT(64'h78887888C0C0C0C0)
) LUT6_2_inst_f0 (
.O6(r[1]),
.O5(r[0]),
.I0(b[1]),
.I1(a[0]),
.I2(b[0]),
.I3(a[1]),
.I4(1'b1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h47777888B8887888)
) LUT6_2_inst_f1 (
.O6(r[2]),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

LUT6_2 #(
.INIT(64'hF8888000C0008000)
) LUT6_2_inst_f2 (
.O6(C1),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

LUT6_2 #(
.INIT(64'h8000000000000000)
) LUT6_2_inst_f3 (
.O6(C0),
.O5(),
.I0(b[2]),
.I1(a[0]),
.I2(b[1]),
.I3(a[1]),
.I4(b[0]),
.I5(a[2]));

/////////STEP0----ORDER0////////////

wire p_s0_o0_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o0_t0_z0_v0 (
.O6(p_s0_o0_0),
.O5(),
.I0(a[3]),
.I1(b[0]),
.I2(a[2]),
.I3(b[1]),
.I4(a[1]),
.I5(b[2]));

wire p_s0_o1_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o0_t0_z1_v0 (
.O6(p_s0_o1_0),
.O5(),
.I0(a[3]),
.I1(b[0]),
.I2(a[2]),
.I3(b[1]),
.I4(a[1]),
.I5(b[2]));

/////////STEP0----ORDER1////////////

/////////STEP0----ORDER2////////////

/////////STEP0----ORDER3////////////

wire p_s0_o3_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o3_t1_z0_v0 (
.O6(p_s0_o3_0),
.O5(),
.I0(a[6]),
.I1(b[0]),
.I2(a[5]),
.I3(b[1]),
.I4(a[4]),
.I5(b[2]));

wire p_s0_o4_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o3_t1_z1_v0 (
.O6(p_s0_o4_0),
.O5(),
.I0(a[6]),
.I1(b[0]),
.I2(a[5]),
.I3(b[1]),
.I4(a[4]),
.I5(b[2]));

/////////STEP0----ORDER4////////////

/////////STEP0----ORDER5////////////

wire p_s0_o5_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o5_t2_z0_v0 (
.O6(p_s0_o5_0),
.O5(),
.I0(a[8]),
.I1(b[0]),
.I2(a[7]),
.I3(b[1]),
.I4(a[6]),
.I5(b[2]));

wire p_s0_o6_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o5_t2_z1_v0 (
.O6(p_s0_o6_0),
.O5(),
.I0(a[8]),
.I1(b[0]),
.I2(a[7]),
.I3(b[1]),
.I4(a[6]),
.I5(b[2]));

/////////STEP0----ORDER6////////////

wire p_s0_o6_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o6_t3_z0_v0 (
.O6(p_s0_o6_1),
.O5(),
.I0(a[9]),
.I1(b[0]),
.I2(a[8]),
.I3(b[1]),
.I4(a[7]),
.I5(b[2]));

wire p_s0_o7_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o6_t3_z1_v0 (
.O6(p_s0_o7_0),
.O5(),
.I0(a[9]),
.I1(b[0]),
.I2(a[8]),
.I3(b[1]),
.I4(a[7]),
.I5(b[2]));

/////////STEP0----ORDER7////////////

/////////STEP0----ORDER8////////////

wire p_s0_o8_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o8_t4_z0_v0 (
.O6(p_s0_o8_0),
.O5(),
.I0(a[11]),
.I1(b[0]),
.I2(a[10]),
.I3(b[1]),
.I4(a[9]),
.I5(b[2]));

wire p_s0_o9_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o8_t4_z1_v0 (
.O6(p_s0_o9_0),
.O5(),
.I0(a[11]),
.I1(b[0]),
.I2(a[10]),
.I3(b[1]),
.I4(a[9]),
.I5(b[2]));

wire p_s0_o8_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o8_t4_z0_v1 (
.O6(p_s0_o8_1),
.O5(),
.I0(a[8]),
.I1(b[3]),
.I2(a[7]),
.I3(b[4]),
.I4(a[6]),
.I5(b[5]));

wire p_s0_o9_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o8_t4_z1_v1 (
.O6(p_s0_o9_1),
.O5(),
.I0(a[8]),
.I1(b[3]),
.I2(a[7]),
.I3(b[4]),
.I4(a[6]),
.I5(b[5]));

/////////STEP0----ORDER9////////////

wire p_s0_o9_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o9_t5_z0_v0 (
.O6(p_s0_o9_2),
.O5(),
.I0(a[12]),
.I1(b[0]),
.I2(a[11]),
.I3(b[1]),
.I4(a[10]),
.I5(b[2]));

wire p_s0_o10_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o9_t5_z1_v0 (
.O6(p_s0_o10_0),
.O5(),
.I0(a[12]),
.I1(b[0]),
.I2(a[11]),
.I3(b[1]),
.I4(a[10]),
.I5(b[2]));

wire p_s0_o9_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o9_t5_z0_v1 (
.O6(p_s0_o9_3),
.O5(),
.I0(a[9]),
.I1(b[3]),
.I2(a[8]),
.I3(b[4]),
.I4(a[7]),
.I5(b[5]));

wire p_s0_o10_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o9_t5_z1_v1 (
.O6(p_s0_o10_1),
.O5(),
.I0(a[9]),
.I1(b[3]),
.I2(a[8]),
.I3(b[4]),
.I4(a[7]),
.I5(b[5]));

/////////STEP0----ORDER10////////////

/////////STEP0----ORDER11////////////

wire p_s0_o11_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o11_t6_z0_v0 (
.O6(p_s0_o11_0),
.O5(),
.I0(a[14]),
.I1(b[0]),
.I2(a[13]),
.I3(b[1]),
.I4(a[12]),
.I5(b[2]));

wire p_s0_o12_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o11_t6_z1_v0 (
.O6(p_s0_o12_0),
.O5(),
.I0(a[14]),
.I1(b[0]),
.I2(a[13]),
.I3(b[1]),
.I4(a[12]),
.I5(b[2]));

wire p_s0_o11_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o11_t6_z0_v1 (
.O6(p_s0_o11_1),
.O5(),
.I0(a[11]),
.I1(b[3]),
.I2(a[10]),
.I3(b[4]),
.I4(a[9]),
.I5(b[5]));

wire p_s0_o12_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o11_t6_z1_v1 (
.O6(p_s0_o12_1),
.O5(),
.I0(a[11]),
.I1(b[3]),
.I2(a[10]),
.I3(b[4]),
.I4(a[9]),
.I5(b[5]));

/////////STEP0----ORDER12////////////

wire p_s0_o12_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o12_t7_z0_v0 (
.O6(p_s0_o12_2),
.O5(),
.I0(a[15]),
.I1(b[0]),
.I2(a[14]),
.I3(b[1]),
.I4(a[13]),
.I5(b[2]));

wire p_s0_o13_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o12_t7_z1_v0 (
.O6(p_s0_o13_0),
.O5(),
.I0(a[15]),
.I1(b[0]),
.I2(a[14]),
.I3(b[1]),
.I4(a[13]),
.I5(b[2]));

wire p_s0_o12_3;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o12_t7_z0_v1 (
.O6(p_s0_o12_3),
.O5(),
.I0(a[12]),
.I1(b[3]),
.I2(a[11]),
.I3(b[4]),
.I4(a[10]),
.I5(b[5]));

wire p_s0_o13_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o12_t7_z1_v1 (
.O6(p_s0_o13_1),
.O5(),
.I0(a[12]),
.I1(b[3]),
.I2(a[11]),
.I3(b[4]),
.I4(a[10]),
.I5(b[5]));

/////////STEP0----ORDER13////////////

wire p_s0_o13_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o13_t8_z0_v0 (
.O6(p_s0_o13_2),
.O5(),
.I0(a[15]),
.I1(b[1]),
.I2(a[14]),
.I3(b[2]),
.I4(a[13]),
.I5(b[3]));

wire p_s0_o14_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o13_t8_z1_v0 (
.O6(p_s0_o14_0),
.O5(),
.I0(a[15]),
.I1(b[1]),
.I2(a[14]),
.I3(b[2]),
.I4(a[13]),
.I5(b[3]));

/////////STEP0----ORDER14////////////

wire p_s0_o14_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o14_t9_z0_v0 (
.O6(p_s0_o14_1),
.O5(),
.I0(a[15]),
.I1(b[2]),
.I2(a[14]),
.I3(b[3]),
.I4(a[13]),
.I5(b[4]));

wire p_s0_o15_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o14_t9_z1_v0 (
.O6(p_s0_o15_0),
.O5(),
.I0(a[15]),
.I1(b[2]),
.I2(a[14]),
.I3(b[3]),
.I4(a[13]),
.I5(b[4]));

wire p_s0_o14_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o14_t9_z0_v1 (
.O6(p_s0_o14_2),
.O5(),
.I0(a[12]),
.I1(b[5]),
.I2(a[11]),
.I3(b[6]),
.I4(a[10]),
.I5(b[7]));

wire p_s0_o15_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o14_t9_z1_v1 (
.O6(p_s0_o15_1),
.O5(),
.I0(a[12]),
.I1(b[5]),
.I2(a[11]),
.I3(b[6]),
.I4(a[10]),
.I5(b[7]));

/////////STEP0----ORDER15////////////

wire p_s0_o15_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o15_t10_z0_v0 (
.O6(p_s0_o15_2),
.O5(),
.I0(a[15]),
.I1(b[3]),
.I2(a[14]),
.I3(b[4]),
.I4(a[13]),
.I5(b[5]));

wire p_s0_o16_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o15_t10_z1_v0 (
.O6(p_s0_o16_0),
.O5(),
.I0(a[15]),
.I1(b[3]),
.I2(a[14]),
.I3(b[4]),
.I4(a[13]),
.I5(b[5]));

/////////STEP0----ORDER16////////////

wire p_s0_o16_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o16_t11_z0_v0 (
.O6(p_s0_o16_1),
.O5(),
.I0(a[15]),
.I1(b[4]),
.I2(a[14]),
.I3(b[5]),
.I4(a[13]),
.I5(b[6]));

wire p_s0_o17_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o16_t11_z1_v0 (
.O6(p_s0_o17_0),
.O5(),
.I0(a[15]),
.I1(b[4]),
.I2(a[14]),
.I3(b[5]),
.I4(a[13]),
.I5(b[6]));

wire p_s0_o16_2;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o16_t11_z0_v1 (
.O6(p_s0_o16_2),
.O5(),
.I0(a[12]),
.I1(b[7]),
.I2(a[11]),
.I3(b[8]),
.I4(a[10]),
.I5(b[9]));

wire p_s0_o17_1;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o16_t11_z1_v1 (
.O6(p_s0_o17_1),
.O5(),
.I0(a[12]),
.I1(b[7]),
.I2(a[11]),
.I3(b[8]),
.I4(a[10]),
.I5(b[9]));

/////////STEP0----ORDER17////////////

/////////STEP0----ORDER18////////////

wire p_s0_o18_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o18_t12_z0_v0 (
.O6(p_s0_o18_0),
.O5(),
.I0(a[15]),
.I1(b[6]),
.I2(a[14]),
.I3(b[7]),
.I4(a[13]),
.I5(b[8]));

wire p_s0_o19_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o18_t12_z1_v0 (
.O6(p_s0_o19_0),
.O5(),
.I0(a[15]),
.I1(b[6]),
.I2(a[14]),
.I3(b[7]),
.I4(a[13]),
.I5(b[8]));

/////////STEP0----ORDER19////////////

wire p_s0_o19_1;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o19_t13_z0_v0 (
.O6(p_s0_o19_1),
.O5(),
.I0(a[15]),
.I1(b[7]),
.I2(a[14]),
.I3(b[8]),
.I4(a[13]),
.I5(b[9]));

wire p_s0_o20_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o19_t13_z1_v0 (
.O6(p_s0_o20_0),
.O5(),
.I0(a[15]),
.I1(b[7]),
.I2(a[14]),
.I3(b[8]),
.I4(a[13]),
.I5(b[9]));

/////////STEP0----ORDER20////////////

/////////STEP0----ORDER21////////////

/////////STEP0----ORDER22////////////

wire p_s0_o22_0;
LUT6_2 #(
.INIT(64'h8777788878887888)
) LUT6_2_inst_s0_o22_t14_z0_v0 (
.O6(p_s0_o22_0),
.O5(),
.I0(a[15]),
.I1(b[10]),
.I2(a[14]),
.I3(b[11]),
.I4(a[13]),
.I5(b[12]));

wire p_s0_o23_0;
LUT6_2 #(
.INIT(64'hF888800080008000)
) LUT6_2_inst_s0_o22_t14_z1_v0 (
.O6(p_s0_o23_0),
.O5(),
.I0(a[15]),
.I1(b[10]),
.I2(a[14]),
.I3(b[11]),
.I4(a[13]),
.I5(b[12]));

/////////STEP0----ORDER23////////////

/////////STEP0----ORDER24////////////

/////////STEP0----ORDER25////////////

/////////STEP0----ORDER26////////////

/////////STEP0----ORDER27////////////

/////////STEP1----ORDER0////////////

/////////STEP1----ORDER1////////////

wire p_s1_o2_0;
wire p_s1_o1_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o1_t15_z0_v0 (
.O6(p_s1_o2_0),
.O5(p_s1_o1_0),
.I0(a[4]),
.I1(b[0]),
.I2(a[3]),
.I3(b[1]),
.I4(p_s0_o1_0),
.I5(1'b1));

/////////STEP1----ORDER2////////////

/////////STEP1----ORDER3////////////

wire p_s1_o4_0;
wire p_s1_o3_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o3_t16_z0_v0 (
.O6(p_s1_o4_0),
.O5(p_s1_o3_0),
.I0(a[3]),
.I1(b[3]),
.I2(a[2]),
.I3(b[4]),
.I4(p_s0_o3_0),
.I5(1'b1));

/////////STEP1----ORDER4////////////

wire p_s1_o5_0;
wire p_s1_o4_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o4_t17_z0_v0 (
.O6(p_s1_o5_0),
.O5(p_s1_o4_1),
.I0(a[7]),
.I1(b[0]),
.I2(a[6]),
.I3(b[1]),
.I4(p_s0_o4_0),
.I5(1'b1));

/////////STEP1----ORDER5////////////

wire p_s1_o6_0;
wire p_s1_o5_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o5_t18_z0_v0 (
.O6(p_s1_o6_0),
.O5(p_s1_o5_1),
.I0(a[5]),
.I1(b[3]),
.I2(a[4]),
.I3(b[4]),
.I4(p_s0_o5_0),
.I5(1'b1));

/////////STEP1----ORDER6////////////

wire p_s1_o7_0;
wire p_s1_o6_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o6_t19_z0_v0 (
.O6(p_s1_o7_0),
.O5(p_s1_o6_1),
.I0(a[6]),
.I1(b[3]),
.I2(a[5]),
.I3(b[4]),
.I4(p_s0_o6_0),
.I5(1'b1));

wire p_s1_o7_1;
wire p_s1_o6_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o6_t19_z0_v1 (
.O6(p_s1_o7_1),
.O5(p_s1_o6_2),
.I0(a[4]),
.I1(b[5]),
.I2(a[3]),
.I3(b[6]),
.I4(p_s0_o6_1),
.I5(1'b1));

/////////STEP1----ORDER7////////////

wire p_s1_o8_0;
wire p_s1_o7_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o7_t20_z0_v0 (
.O6(p_s1_o8_0),
.O5(p_s1_o7_2),
.I0(a[10]),
.I1(b[0]),
.I2(a[9]),
.I3(b[1]),
.I4(p_s0_o7_0),
.I5(1'b1));

/////////STEP1----ORDER8////////////

wire p_s1_o9_0;
wire p_s1_o8_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o8_t21_z0_v0 (
.O6(p_s1_o9_0),
.O5(p_s1_o8_1),
.I0(a[5]),
.I1(b[6]),
.I2(a[4]),
.I3(b[7]),
.I4(p_s0_o8_0),
.I5(1'b1));

/////////STEP1----ORDER9////////////

wire p_s1_o10_0;
wire p_s1_o9_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o9_t22_z0_v0 (
.O6(p_s1_o10_0),
.O5(p_s1_o9_1),
.I0(a[6]),
.I1(b[6]),
.I2(a[5]),
.I3(b[7]),
.I4(p_s0_o9_0),
.I5(1'b1));

wire p_s1_o10_1;
wire p_s1_o9_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o9_t22_z0_v1 (
.O6(p_s1_o10_1),
.O5(p_s1_o9_2),
.I0(a[4]),
.I1(b[8]),
.I2(a[3]),
.I3(b[9]),
.I4(p_s0_o9_1),
.I5(1'b1));

wire p_s1_o10_2;
wire p_s1_o9_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o9_t22_z0_v2 (
.O6(p_s1_o10_2),
.O5(p_s1_o9_3),
.I0(a[2]),
.I1(b[10]),
.I2(a[1]),
.I3(b[11]),
.I4(p_s0_o9_2),
.I5(1'b1));

/////////STEP1----ORDER10////////////

wire p_s1_o11_0;
wire p_s1_o10_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o10_t23_z0_v0 (
.O6(p_s1_o11_0),
.O5(p_s1_o10_3),
.I0(a[13]),
.I1(b[0]),
.I2(a[12]),
.I3(b[1]),
.I4(p_s0_o10_0),
.I5(1'b1));

wire p_s1_o11_1;
wire p_s1_o10_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o10_t23_z0_v1 (
.O6(p_s1_o11_1),
.O5(p_s1_o10_4),
.I0(a[11]),
.I1(b[2]),
.I2(a[10]),
.I3(b[3]),
.I4(p_s0_o10_1),
.I5(1'b1));

/////////STEP1----ORDER11////////////

wire p_s1_o12_0;
wire p_s1_o11_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o11_t24_z0_v0 (
.O6(p_s1_o12_0),
.O5(p_s1_o11_2),
.I0(a[8]),
.I1(b[6]),
.I2(a[7]),
.I3(b[7]),
.I4(p_s0_o11_0),
.I5(1'b1));

wire p_s1_o12_1;
wire p_s1_o11_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o11_t24_z0_v1 (
.O6(p_s1_o12_1),
.O5(p_s1_o11_3),
.I0(a[6]),
.I1(b[8]),
.I2(a[5]),
.I3(b[9]),
.I4(p_s0_o11_1),
.I5(1'b1));

/////////STEP1----ORDER12////////////

wire p_s1_o13_0;
wire p_s1_o12_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o12_t25_z0_v0 (
.O6(p_s1_o13_0),
.O5(p_s1_o12_2),
.I0(a[9]),
.I1(b[6]),
.I2(a[8]),
.I3(b[7]),
.I4(p_s0_o12_0),
.I5(1'b1));

wire p_s1_o13_1;
wire p_s1_o12_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o12_t25_z0_v1 (
.O6(p_s1_o13_1),
.O5(p_s1_o12_3),
.I0(a[7]),
.I1(b[8]),
.I2(a[6]),
.I3(b[9]),
.I4(p_s0_o12_1),
.I5(1'b1));

wire p_s1_o13_2;
wire p_s1_o12_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o12_t25_z0_v2 (
.O6(p_s1_o13_2),
.O5(p_s1_o12_4),
.I0(a[5]),
.I1(b[10]),
.I2(a[4]),
.I3(b[11]),
.I4(p_s0_o12_2),
.I5(1'b1));

wire p_s1_o13_3;
wire p_s1_o12_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o12_t25_z0_v3 (
.O6(p_s1_o13_3),
.O5(p_s1_o12_5),
.I0(a[3]),
.I1(b[12]),
.I2(a[2]),
.I3(b[13]),
.I4(p_s0_o12_3),
.I5(1'b1));

/////////STEP1----ORDER13////////////

wire p_s1_o14_0;
wire p_s1_o13_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o13_t26_z0_v0 (
.O6(p_s1_o14_0),
.O5(p_s1_o13_4),
.I0(a[12]),
.I1(b[4]),
.I2(a[11]),
.I3(b[5]),
.I4(p_s0_o13_0),
.I5(1'b1));

wire p_s1_o14_1;
wire p_s1_o13_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o13_t26_z0_v1 (
.O6(p_s1_o14_1),
.O5(p_s1_o13_5),
.I0(a[10]),
.I1(b[6]),
.I2(a[9]),
.I3(b[7]),
.I4(p_s0_o13_1),
.I5(1'b1));

wire p_s1_o14_2;
wire p_s1_o13_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o13_t26_z0_v2 (
.O6(p_s1_o14_2),
.O5(p_s1_o13_6),
.I0(a[8]),
.I1(b[8]),
.I2(a[7]),
.I3(b[9]),
.I4(p_s0_o13_2),
.I5(1'b1));

/////////STEP1----ORDER14////////////

wire p_s1_o15_0;
wire p_s1_o14_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t27_z0_v0 (
.O6(p_s1_o15_0),
.O5(p_s1_o14_3),
.I0(a[9]),
.I1(b[8]),
.I2(a[8]),
.I3(b[9]),
.I4(p_s0_o14_0),
.I5(1'b1));

wire p_s1_o15_1;
wire p_s1_o14_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t27_z0_v1 (
.O6(p_s1_o15_1),
.O5(p_s1_o14_4),
.I0(a[7]),
.I1(b[10]),
.I2(a[6]),
.I3(b[11]),
.I4(p_s0_o14_1),
.I5(1'b1));

wire p_s1_o15_2;
wire p_s1_o14_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o14_t27_z0_v2 (
.O6(p_s1_o15_2),
.O5(p_s1_o14_5),
.I0(a[5]),
.I1(b[12]),
.I2(a[4]),
.I3(b[13]),
.I4(p_s0_o14_2),
.I5(1'b1));

/////////STEP1----ORDER15////////////

wire p_s1_o16_0;
wire p_s1_o15_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o15_t28_z0_v0 (
.O6(p_s1_o16_0),
.O5(p_s1_o15_3),
.I0(a[12]),
.I1(b[6]),
.I2(a[11]),
.I3(b[7]),
.I4(p_s0_o15_0),
.I5(1'b1));

wire p_s1_o16_1;
wire p_s1_o15_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o15_t28_z0_v1 (
.O6(p_s1_o16_1),
.O5(p_s1_o15_4),
.I0(a[10]),
.I1(b[8]),
.I2(a[9]),
.I3(b[9]),
.I4(p_s0_o15_1),
.I5(1'b1));

wire p_s1_o16_2;
wire p_s1_o15_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o15_t28_z0_v2 (
.O6(p_s1_o16_2),
.O5(p_s1_o15_5),
.I0(a[8]),
.I1(b[10]),
.I2(a[7]),
.I3(b[11]),
.I4(p_s0_o15_2),
.I5(1'b1));

/////////STEP1----ORDER16////////////

wire p_s1_o17_0;
wire p_s1_o16_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o16_t29_z0_v0 (
.O6(p_s1_o17_0),
.O5(p_s1_o16_3),
.I0(a[9]),
.I1(b[10]),
.I2(a[8]),
.I3(b[11]),
.I4(p_s0_o16_0),
.I5(1'b1));

wire p_s1_o17_1;
wire p_s1_o16_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o16_t29_z0_v1 (
.O6(p_s1_o17_1),
.O5(p_s1_o16_4),
.I0(a[7]),
.I1(b[12]),
.I2(a[6]),
.I3(b[13]),
.I4(p_s0_o16_1),
.I5(1'b1));

wire p_s1_o17_2;
wire p_s1_o16_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o16_t29_z0_v2 (
.O6(p_s1_o17_2),
.O5(p_s1_o16_5),
.I0(a[5]),
.I1(b[14]),
.I2(a[4]),
.I3(b[15]),
.I4(p_s0_o16_2),
.I5(1'b1));

/////////STEP1----ORDER17////////////

wire p_s1_o18_0;
wire p_s1_o17_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o17_t30_z0_v0 (
.O6(p_s1_o18_0),
.O5(p_s1_o17_3),
.I0(a[15]),
.I1(b[5]),
.I2(a[14]),
.I3(b[6]),
.I4(p_s0_o17_0),
.I5(1'b1));

wire p_s1_o18_1;
wire p_s1_o17_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o17_t30_z0_v1 (
.O6(p_s1_o18_1),
.O5(p_s1_o17_4),
.I0(a[13]),
.I1(b[7]),
.I2(a[12]),
.I3(b[8]),
.I4(p_s0_o17_1),
.I5(1'b1));

/////////STEP1----ORDER18////////////

wire p_s1_o19_0;
wire p_s1_o18_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o18_t31_z0_v0 (
.O6(p_s1_o19_0),
.O5(p_s1_o18_2),
.I0(a[12]),
.I1(b[9]),
.I2(a[11]),
.I3(b[10]),
.I4(p_s0_o18_0),
.I5(1'b1));

/////////STEP1----ORDER19////////////

wire p_s1_o20_0;
wire p_s1_o19_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t32_z0_v0 (
.O6(p_s1_o20_0),
.O5(p_s1_o19_1),
.I0(a[12]),
.I1(b[10]),
.I2(a[11]),
.I3(b[11]),
.I4(p_s0_o19_0),
.I5(1'b1));

wire p_s1_o20_1;
wire p_s1_o19_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o19_t32_z0_v1 (
.O6(p_s1_o20_1),
.O5(p_s1_o19_2),
.I0(a[10]),
.I1(b[12]),
.I2(a[9]),
.I3(b[13]),
.I4(p_s0_o19_1),
.I5(1'b1));

/////////STEP1----ORDER20////////////

wire p_s1_o21_0;
wire p_s1_o20_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o20_t33_z0_v0 (
.O6(p_s1_o21_0),
.O5(p_s1_o20_2),
.I0(a[15]),
.I1(b[8]),
.I2(a[14]),
.I3(b[9]),
.I4(p_s0_o20_0),
.I5(1'b1));

/////////STEP1----ORDER21////////////

/////////STEP1----ORDER22////////////

wire p_s1_o23_0;
wire p_s1_o22_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o22_t34_z0_v0 (
.O6(p_s1_o23_0),
.O5(p_s1_o22_0),
.I0(a[12]),
.I1(b[13]),
.I2(a[11]),
.I3(b[14]),
.I4(p_s0_o22_0),
.I5(1'b1));

/////////STEP1----ORDER23////////////

wire p_s1_o24_0;
wire p_s1_o23_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s1_o23_t35_z0_v0 (
.O6(p_s1_o24_0),
.O5(p_s1_o23_1),
.I0(a[15]),
.I1(b[11]),
.I2(a[14]),
.I3(b[12]),
.I4(p_s0_o23_0),
.I5(1'b1));

/////////STEP1----ORDER24////////////

/////////STEP1----ORDER25////////////

/////////STEP1----ORDER26////////////

/////////STEP1----ORDER27////////////

/////////STEP2----ORDER0////////////

/////////STEP2----ORDER1////////////

wire p_s2_o2_0;
wire p_s2_o1_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o1_t43_z0_v0 (
.O6(p_s2_o2_0),
.O5(p_s2_o1_0),
.I0(a[2]),
.I1(b[2]),
.I2(a[1]),
.I3(b[3]),
.I4(p_s1_o1_0),
.I5(1'b1));

/////////STEP2----ORDER2////////////

wire p_s2_o3_0;
wire p_s2_o2_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o2_t44_z0_v0 (
.O6(p_s2_o3_0),
.O5(p_s2_o2_1),
.I0(a[5]),
.I1(b[0]),
.I2(a[4]),
.I3(b[1]),
.I4(p_s1_o2_0),
.I5(1'b1));

/////////STEP2----ORDER3////////////

wire p_s2_o4_0;
wire p_s2_o3_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o3_t45_z0_v0 (
.O6(p_s2_o4_0),
.O5(p_s2_o3_1),
.I0(a[1]),
.I1(b[5]),
.I2(a[0]),
.I3(b[6]),
.I4(p_s1_o3_0),
.I5(1'b1));

/////////STEP2----ORDER4////////////

wire p_s2_o5_0;
wire p_s2_o4_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o4_t46_z0_v0 (
.O6(p_s2_o5_0),
.O5(p_s2_o4_1),
.I0(a[5]),
.I1(b[2]),
.I2(a[4]),
.I3(b[3]),
.I4(p_s1_o4_0),
.I5(1'b1));

wire p_s2_o5_1;
wire p_s2_o4_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o4_t46_z0_v1 (
.O6(p_s2_o5_1),
.O5(p_s2_o4_2),
.I0(a[3]),
.I1(b[4]),
.I2(a[2]),
.I3(b[5]),
.I4(p_s1_o4_1),
.I5(1'b1));

/////////STEP2----ORDER5////////////

wire p_s2_o6_0;
wire p_s2_o5_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o5_t47_z0_v0 (
.O6(p_s2_o6_0),
.O5(p_s2_o5_2),
.I0(a[3]),
.I1(b[5]),
.I2(a[2]),
.I3(b[6]),
.I4(p_s1_o5_0),
.I5(1'b1));

wire p_s2_o6_1;
wire p_s2_o5_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o5_t47_z0_v1 (
.O6(p_s2_o6_1),
.O5(p_s2_o5_3),
.I0(a[1]),
.I1(b[7]),
.I2(a[0]),
.I3(b[8]),
.I4(p_s1_o5_1),
.I5(1'b1));

/////////STEP2----ORDER6////////////

wire p_s2_o7_0;
wire p_s2_o6_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o6_t48_z0_v0 (
.O6(p_s2_o7_0),
.O5(p_s2_o6_2),
.I0(a[2]),
.I1(b[7]),
.I2(a[1]),
.I3(b[8]),
.I4(p_s1_o6_0),
.I5(1'b1));

/////////STEP2----ORDER7////////////

wire p_s2_o8_0;
wire p_s2_o7_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o7_t49_z0_v0 (
.O6(p_s2_o8_0),
.O5(p_s2_o7_1),
.I0(a[8]),
.I1(b[2]),
.I2(a[7]),
.I3(b[3]),
.I4(p_s1_o7_0),
.I5(1'b1));

wire p_s2_o8_1;
wire p_s2_o7_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o7_t49_z0_v1 (
.O6(p_s2_o8_1),
.O5(p_s2_o7_2),
.I0(a[6]),
.I1(b[4]),
.I2(a[5]),
.I3(b[5]),
.I4(p_s1_o7_1),
.I5(1'b1));

wire p_s2_o8_2;
wire p_s2_o7_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o7_t49_z0_v2 (
.O6(p_s2_o8_2),
.O5(p_s2_o7_3),
.I0(a[4]),
.I1(b[6]),
.I2(a[3]),
.I3(b[7]),
.I4(p_s1_o7_2),
.I5(1'b1));

/////////STEP2----ORDER8////////////

wire p_s2_o9_0;
wire p_s2_o8_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o8_t50_z0_v0 (
.O6(p_s2_o9_0),
.O5(p_s2_o8_3),
.I0(a[3]),
.I1(b[8]),
.I2(a[2]),
.I3(b[9]),
.I4(p_s1_o8_0),
.I5(1'b1));

wire p_s2_o9_1;
wire p_s2_o8_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o8_t50_z0_v1 (
.O6(p_s2_o9_1),
.O5(p_s2_o8_4),
.I0(a[1]),
.I1(b[10]),
.I2(a[0]),
.I3(b[11]),
.I4(p_s1_o8_1),
.I5(1'b1));

/////////STEP2----ORDER9////////////

wire p_s2_o10_0;
wire p_s2_o9_2;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o9_t39_z0_v0 (
.O6(p_s2_o10_0),
.O5(p_s2_o9_2),
.I0(a[0]),
.I1(b[12]),
.I2(p_s1_o9_0),
.I3(p_s1_o9_1),
.I4(1'b0),
.I5(1'b1));

/////////STEP2----ORDER10////////////

wire p_s2_o11_0;
wire p_s2_o10_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o10_t51_z0_v0 (
.O6(p_s2_o11_0),
.O5(p_s2_o10_1),
.I0(a[9]),
.I1(b[4]),
.I2(a[8]),
.I3(b[5]),
.I4(p_s1_o10_0),
.I5(1'b1));

wire p_s2_o11_1;
wire p_s2_o10_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o10_t51_z0_v1 (
.O6(p_s2_o11_1),
.O5(p_s2_o10_2),
.I0(a[7]),
.I1(b[6]),
.I2(a[6]),
.I3(b[7]),
.I4(p_s1_o10_1),
.I5(1'b1));

wire p_s2_o11_2;
wire p_s2_o10_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o10_t51_z0_v2 (
.O6(p_s2_o11_2),
.O5(p_s2_o10_3),
.I0(a[5]),
.I1(b[8]),
.I2(a[4]),
.I3(b[9]),
.I4(p_s1_o10_2),
.I5(1'b1));

wire p_s2_o11_3;
wire p_s2_o10_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o10_t51_z0_v3 (
.O6(p_s2_o11_3),
.O5(p_s2_o10_4),
.I0(a[3]),
.I1(b[10]),
.I2(a[2]),
.I3(b[11]),
.I4(p_s1_o10_3),
.I5(1'b1));

wire p_s2_o11_4;
wire p_s2_o10_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o10_t51_z0_v4 (
.O6(p_s2_o11_4),
.O5(p_s2_o10_5),
.I0(a[1]),
.I1(b[12]),
.I2(a[0]),
.I3(b[13]),
.I4(p_s1_o10_4),
.I5(1'b1));

/////////STEP2----ORDER11////////////

wire p_s2_o12_0;
wire p_s2_o11_5;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o11_t40_z0_v0 (
.O6(p_s2_o12_0),
.O5(p_s2_o11_5),
.I0(a[4]),
.I1(b[10]),
.I2(p_s1_o11_0),
.I3(p_s1_o11_1),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o12_1;
wire p_s2_o11_6;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o11_t52_z0_v0 (
.O6(p_s2_o12_1),
.O5(p_s2_o11_6),
.I0(a[3]),
.I1(b[11]),
.I2(a[2]),
.I3(b[12]),
.I4(p_s1_o11_2),
.I5(1'b1));

wire p_s2_o12_2;
wire p_s2_o11_7;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o11_t52_z0_v1 (
.O6(p_s2_o12_2),
.O5(p_s2_o11_7),
.I0(a[1]),
.I1(b[13]),
.I2(a[0]),
.I3(b[14]),
.I4(p_s1_o11_3),
.I5(1'b1));

/////////STEP2----ORDER12////////////

wire p_s2_o13_0;
wire p_s2_o12_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o12_t53_z0_v0 (
.O6(p_s2_o13_0),
.O5(p_s2_o12_3),
.I0(a[1]),
.I1(b[14]),
.I2(a[0]),
.I3(b[15]),
.I4(p_s1_o12_0),
.I5(1'b1));

wire p_s2_o12_4;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o12_t64_z0_v0 (
.O6(p_s2_o12_4),
.O5(),
.I0(p_s1_o12_1),
.I1(p_s1_o12_2),
.I2(p_s1_o12_3),
.I3(p_s1_o12_4),
.I4(p_s1_o12_5),
.I5(p_s1_o13_0));

wire p_s2_o13_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o12_t64_z1_v0 (
.O6(p_s2_o13_1),
.O5(),
.I0(p_s1_o12_1),
.I1(p_s1_o12_2),
.I2(p_s1_o12_3),
.I3(p_s1_o12_4),
.I4(p_s1_o12_5),
.I5(p_s1_o13_0));

wire p_s2_o14_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o12_t64_z2_v0 (
.O6(p_s2_o14_0),
.O5(),
.I0(p_s1_o12_1),
.I1(p_s1_o12_2),
.I2(p_s1_o12_3),
.I3(p_s1_o12_4),
.I4(p_s1_o12_5),
.I5(p_s1_o13_0));

/////////STEP2----ORDER13////////////

wire p_s2_o14_1;
wire p_s2_o13_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s2_o13_t36_z0_v0 (
.O6(p_s2_o14_1),
.O5(p_s2_o13_2),
.I0(p_s1_o13_1),
.I1(p_s1_o13_2),
.I2(p_s1_o13_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o14_2;
wire p_s2_o13_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o13_t54_z0_v0 (
.O6(p_s2_o14_2),
.O5(p_s2_o13_3),
.I0(a[6]),
.I1(b[10]),
.I2(a[5]),
.I3(b[11]),
.I4(p_s1_o13_4),
.I5(1'b1));

wire p_s2_o14_3;
wire p_s2_o13_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o13_t54_z0_v1 (
.O6(p_s2_o14_3),
.O5(p_s2_o13_4),
.I0(a[4]),
.I1(b[12]),
.I2(a[3]),
.I3(b[13]),
.I4(p_s1_o13_5),
.I5(1'b1));

wire p_s2_o14_4;
wire p_s2_o13_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o13_t54_z0_v2 (
.O6(p_s2_o14_4),
.O5(p_s2_o13_5),
.I0(a[2]),
.I1(b[14]),
.I2(a[1]),
.I3(b[15]),
.I4(p_s1_o13_6),
.I5(1'b1));

/////////STEP2----ORDER14////////////

wire p_s2_o15_0;
wire p_s2_o14_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o14_t55_z0_v0 (
.O6(p_s2_o15_0),
.O5(p_s2_o14_5),
.I0(a[3]),
.I1(b[14]),
.I2(a[2]),
.I3(b[15]),
.I4(p_s1_o14_0),
.I5(1'b1));

wire p_s2_o14_6;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s2_o14_t65_z0_v0 (
.O6(p_s2_o14_6),
.O5(),
.I0(p_s1_o14_1),
.I1(p_s1_o14_2),
.I2(p_s1_o14_3),
.I3(p_s1_o14_4),
.I4(p_s1_o14_5),
.I5(p_s1_o15_0));

wire p_s2_o15_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s2_o14_t65_z1_v0 (
.O6(p_s2_o15_1),
.O5(),
.I0(p_s1_o14_1),
.I1(p_s1_o14_2),
.I2(p_s1_o14_3),
.I3(p_s1_o14_4),
.I4(p_s1_o14_5),
.I5(p_s1_o15_0));

wire p_s2_o16_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s2_o14_t65_z2_v0 (
.O6(p_s2_o16_0),
.O5(),
.I0(p_s1_o14_1),
.I1(p_s1_o14_2),
.I2(p_s1_o14_3),
.I3(p_s1_o14_4),
.I4(p_s1_o14_5),
.I5(p_s1_o15_0));

/////////STEP2----ORDER15////////////

wire p_s2_o16_1;
wire p_s2_o15_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s2_o15_t37_z0_v0 (
.O6(p_s2_o16_1),
.O5(p_s2_o15_2),
.I0(p_s1_o15_1),
.I1(p_s1_o15_2),
.I2(p_s1_o15_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o16_2;
wire p_s2_o15_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o15_t56_z0_v0 (
.O6(p_s2_o16_2),
.O5(p_s2_o15_3),
.I0(a[6]),
.I1(b[12]),
.I2(a[5]),
.I3(b[13]),
.I4(p_s1_o15_4),
.I5(1'b1));

wire p_s2_o16_3;
wire p_s2_o15_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o15_t56_z0_v1 (
.O6(p_s2_o16_3),
.O5(p_s2_o15_4),
.I0(a[4]),
.I1(b[14]),
.I2(a[3]),
.I3(b[15]),
.I4(p_s1_o15_5),
.I5(1'b1));

/////////STEP2----ORDER16////////////

wire p_s2_o17_0;
wire p_s2_o16_4;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s2_o16_t38_z0_v0 (
.O6(p_s2_o17_0),
.O5(p_s2_o16_4),
.I0(p_s1_o16_0),
.I1(p_s1_o16_1),
.I2(p_s1_o16_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o17_1;
wire p_s2_o16_5;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s2_o16_t38_z0_v1 (
.O6(p_s2_o17_1),
.O5(p_s2_o16_5),
.I0(p_s1_o16_3),
.I1(p_s1_o16_4),
.I2(p_s1_o16_5),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP2----ORDER17////////////

wire p_s2_o18_0;
wire p_s2_o17_2;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o17_t41_z0_v0 (
.O6(p_s2_o18_0),
.O5(p_s2_o17_2),
.I0(a[11]),
.I1(b[9]),
.I2(p_s1_o17_0),
.I3(p_s1_o17_1),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o18_1;
wire p_s2_o17_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o17_t57_z0_v0 (
.O6(p_s2_o18_1),
.O5(p_s2_o17_3),
.I0(a[10]),
.I1(b[10]),
.I2(a[9]),
.I3(b[11]),
.I4(p_s1_o17_2),
.I5(1'b1));

wire p_s2_o18_2;
wire p_s2_o17_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o17_t57_z0_v1 (
.O6(p_s2_o18_2),
.O5(p_s2_o17_4),
.I0(a[8]),
.I1(b[12]),
.I2(a[7]),
.I3(b[13]),
.I4(p_s1_o17_3),
.I5(1'b1));

wire p_s2_o18_3;
wire p_s2_o17_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o17_t57_z0_v2 (
.O6(p_s2_o18_3),
.O5(p_s2_o17_5),
.I0(a[6]),
.I1(b[14]),
.I2(a[5]),
.I3(b[15]),
.I4(p_s1_o17_4),
.I5(1'b1));

/////////STEP2----ORDER18////////////

wire p_s2_o19_0;
wire p_s2_o18_4;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s2_o18_t42_z0_v0 (
.O6(p_s2_o19_0),
.O5(p_s2_o18_4),
.I0(a[10]),
.I1(b[11]),
.I2(p_s1_o18_0),
.I3(p_s1_o18_1),
.I4(1'b0),
.I5(1'b1));

wire p_s2_o19_1;
wire p_s2_o18_5;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o18_t58_z0_v0 (
.O6(p_s2_o19_1),
.O5(p_s2_o18_5),
.I0(a[9]),
.I1(b[12]),
.I2(a[8]),
.I3(b[13]),
.I4(p_s1_o18_2),
.I5(1'b1));

/////////STEP2----ORDER19////////////

wire p_s2_o20_0;
wire p_s2_o19_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o19_t59_z0_v0 (
.O6(p_s2_o20_0),
.O5(p_s2_o19_2),
.I0(a[8]),
.I1(b[14]),
.I2(a[7]),
.I3(b[15]),
.I4(p_s1_o19_0),
.I5(1'b1));

/////////STEP2----ORDER20////////////

wire p_s2_o21_0;
wire p_s2_o20_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o20_t60_z0_v0 (
.O6(p_s2_o21_0),
.O5(p_s2_o20_1),
.I0(a[13]),
.I1(b[10]),
.I2(a[12]),
.I3(b[11]),
.I4(p_s1_o20_0),
.I5(1'b1));

wire p_s2_o21_1;
wire p_s2_o20_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o20_t60_z0_v1 (
.O6(p_s2_o21_1),
.O5(p_s2_o20_2),
.I0(a[11]),
.I1(b[12]),
.I2(a[10]),
.I3(b[13]),
.I4(p_s1_o20_1),
.I5(1'b1));

wire p_s2_o21_2;
wire p_s2_o20_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o20_t60_z0_v2 (
.O6(p_s2_o21_2),
.O5(p_s2_o20_3),
.I0(a[9]),
.I1(b[14]),
.I2(a[8]),
.I3(b[15]),
.I4(p_s1_o20_2),
.I5(1'b1));

/////////STEP2----ORDER21////////////

wire p_s2_o22_0;
wire p_s2_o21_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o21_t61_z0_v0 (
.O6(p_s2_o22_0),
.O5(p_s2_o21_3),
.I0(a[15]),
.I1(b[9]),
.I2(a[14]),
.I3(b[10]),
.I4(p_s1_o21_0),
.I5(1'b1));

/////////STEP2----ORDER22////////////

/////////STEP2----ORDER23////////////

wire p_s2_o24_0;
wire p_s2_o23_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o23_t62_z0_v0 (
.O6(p_s2_o24_0),
.O5(p_s2_o23_0),
.I0(a[13]),
.I1(b[13]),
.I2(a[12]),
.I3(b[14]),
.I4(p_s1_o23_0),
.I5(1'b1));

/////////STEP2----ORDER24////////////

wire p_s2_o25_0;
wire p_s2_o24_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s2_o24_t63_z0_v0 (
.O6(p_s2_o25_0),
.O5(p_s2_o24_1),
.I0(a[15]),
.I1(b[12]),
.I2(a[14]),
.I3(b[13]),
.I4(p_s1_o24_0),
.I5(1'b1));

/////////STEP2----ORDER25////////////

/////////STEP2----ORDER26////////////

/////////STEP2----ORDER27////////////

/////////STEP3----ORDER0////////////

/////////STEP3----ORDER1////////////

/////////STEP3----ORDER2////////////

wire p_s3_o3_0;
wire p_s3_o2_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o2_t74_z0_v0 (
.O6(p_s3_o3_0),
.O5(p_s3_o2_0),
.I0(a[3]),
.I1(b[2]),
.I2(a[2]),
.I3(b[3]),
.I4(p_s2_o2_0),
.I5(1'b1));

wire p_s3_o3_1;
wire p_s3_o2_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o2_t74_z0_v1 (
.O6(p_s3_o3_1),
.O5(p_s3_o2_1),
.I0(a[1]),
.I1(b[4]),
.I2(a[0]),
.I3(b[5]),
.I4(p_s2_o2_1),
.I5(1'b1));

/////////STEP3----ORDER3////////////

/////////STEP3----ORDER4////////////

wire p_s3_o5_0;
wire p_s3_o4_0;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o4_t75_z0_v0 (
.O6(p_s3_o5_0),
.O5(p_s3_o4_0),
.I0(a[1]),
.I1(b[6]),
.I2(a[0]),
.I3(b[7]),
.I4(p_s2_o4_0),
.I5(1'b1));

/////////STEP3----ORDER5////////////

/////////STEP3----ORDER6////////////

wire p_s3_o6_0;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o6_t81_z0_v0 (
.O6(p_s3_o6_0),
.O5(),
.I0(p_s2_o6_0),
.I1(p_s2_o6_1),
.I2(p_s2_o6_2),
.I3(p_s1_o6_1),
.I4(p_s1_o6_2),
.I5(p_s2_o7_0));

wire p_s3_o7_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o6_t81_z1_v0 (
.O6(p_s3_o7_0),
.O5(),
.I0(p_s2_o6_0),
.I1(p_s2_o6_1),
.I2(p_s2_o6_2),
.I3(p_s1_o6_1),
.I4(p_s1_o6_2),
.I5(p_s2_o7_0));

wire p_s3_o8_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o6_t81_z2_v0 (
.O6(p_s3_o8_0),
.O5(),
.I0(p_s2_o6_0),
.I1(p_s2_o6_1),
.I2(p_s2_o6_2),
.I3(p_s1_o6_1),
.I4(p_s1_o6_2),
.I5(p_s2_o7_0));

/////////STEP3----ORDER7////////////

wire p_s3_o8_1;
wire p_s3_o7_1;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o7_t70_z0_v0 (
.O6(p_s3_o8_1),
.O5(p_s3_o7_1),
.I0(a[2]),
.I1(b[8]),
.I2(p_s2_o7_1),
.I3(p_s2_o7_2),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o8_2;
wire p_s3_o7_2;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o7_t76_z0_v0 (
.O6(p_s3_o8_2),
.O5(p_s3_o7_2),
.I0(a[1]),
.I1(b[9]),
.I2(a[0]),
.I3(b[10]),
.I4(p_s2_o7_3),
.I5(1'b1));

/////////STEP3----ORDER8////////////

wire p_s3_o8_3;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o8_t82_z0_v0 (
.O6(p_s3_o8_3),
.O5(),
.I0(p_s2_o8_0),
.I1(p_s2_o8_1),
.I2(p_s2_o8_2),
.I3(p_s2_o8_3),
.I4(p_s2_o8_4),
.I5(p_s2_o9_0));

wire p_s3_o9_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o8_t82_z1_v0 (
.O6(p_s3_o9_0),
.O5(),
.I0(p_s2_o8_0),
.I1(p_s2_o8_1),
.I2(p_s2_o8_2),
.I3(p_s2_o8_3),
.I4(p_s2_o8_4),
.I5(p_s2_o9_0));

wire p_s3_o10_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o8_t82_z2_v0 (
.O6(p_s3_o10_0),
.O5(),
.I0(p_s2_o8_0),
.I1(p_s2_o8_1),
.I2(p_s2_o8_2),
.I3(p_s2_o8_3),
.I4(p_s2_o8_4),
.I5(p_s2_o9_0));

/////////STEP3----ORDER9////////////

wire p_s3_o9_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o9_t83_z0_v0 (
.O6(p_s3_o9_1),
.O5(),
.I0(p_s2_o9_1),
.I1(p_s2_o9_2),
.I2(p_s1_o9_2),
.I3(p_s1_o9_3),
.I4(p_s0_o9_3),
.I5(p_s2_o10_0));

wire p_s3_o10_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o9_t83_z1_v0 (
.O6(p_s3_o10_1),
.O5(),
.I0(p_s2_o9_1),
.I1(p_s2_o9_2),
.I2(p_s1_o9_2),
.I3(p_s1_o9_3),
.I4(p_s0_o9_3),
.I5(p_s2_o10_0));

wire p_s3_o11_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o9_t83_z2_v0 (
.O6(p_s3_o11_0),
.O5(),
.I0(p_s2_o9_1),
.I1(p_s2_o9_2),
.I2(p_s1_o9_2),
.I3(p_s1_o9_3),
.I4(p_s0_o9_3),
.I5(p_s2_o10_0));

/////////STEP3----ORDER10////////////

wire p_s3_o10_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o10_t84_z0_v0 (
.O6(p_s3_o10_2),
.O5(),
.I0(p_s2_o10_1),
.I1(p_s2_o10_2),
.I2(p_s2_o10_3),
.I3(p_s2_o10_4),
.I4(p_s2_o10_5),
.I5(p_s2_o11_0));

wire p_s3_o11_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o10_t84_z1_v0 (
.O6(p_s3_o11_1),
.O5(),
.I0(p_s2_o10_1),
.I1(p_s2_o10_2),
.I2(p_s2_o10_3),
.I3(p_s2_o10_4),
.I4(p_s2_o10_5),
.I5(p_s2_o11_0));

wire p_s3_o12_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o10_t84_z2_v0 (
.O6(p_s3_o12_0),
.O5(),
.I0(p_s2_o10_1),
.I1(p_s2_o10_2),
.I2(p_s2_o10_3),
.I3(p_s2_o10_4),
.I4(p_s2_o10_5),
.I5(p_s2_o11_0));

/////////STEP3----ORDER11////////////

wire p_s3_o12_1;
wire p_s3_o11_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o11_t66_z0_v0 (
.O6(p_s3_o12_1),
.O5(p_s3_o11_2),
.I0(p_s2_o11_1),
.I1(p_s2_o11_2),
.I2(p_s2_o11_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o12_2;
wire p_s3_o11_3;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o11_t66_z0_v1 (
.O6(p_s3_o12_2),
.O5(p_s3_o11_3),
.I0(p_s2_o11_4),
.I1(p_s2_o11_5),
.I2(p_s2_o11_6),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER12////////////

wire p_s3_o12_3;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o12_t85_z0_v0 (
.O6(p_s3_o12_3),
.O5(),
.I0(p_s2_o12_0),
.I1(p_s2_o12_1),
.I2(p_s2_o12_2),
.I3(p_s2_o12_3),
.I4(p_s2_o12_4),
.I5(p_s2_o13_0));

wire p_s3_o13_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o12_t85_z1_v0 (
.O6(p_s3_o13_0),
.O5(),
.I0(p_s2_o12_0),
.I1(p_s2_o12_1),
.I2(p_s2_o12_2),
.I3(p_s2_o12_3),
.I4(p_s2_o12_4),
.I5(p_s2_o13_0));

wire p_s3_o14_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o12_t85_z2_v0 (
.O6(p_s3_o14_0),
.O5(),
.I0(p_s2_o12_0),
.I1(p_s2_o12_1),
.I2(p_s2_o12_2),
.I3(p_s2_o12_3),
.I4(p_s2_o12_4),
.I5(p_s2_o13_0));

/////////STEP3----ORDER13////////////

wire p_s3_o13_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o13_t86_z0_v0 (
.O6(p_s3_o13_1),
.O5(),
.I0(p_s2_o13_1),
.I1(p_s2_o13_2),
.I2(p_s2_o13_3),
.I3(p_s2_o13_4),
.I4(p_s2_o13_5),
.I5(p_s2_o14_0));

wire p_s3_o14_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o13_t86_z1_v0 (
.O6(p_s3_o14_1),
.O5(),
.I0(p_s2_o13_1),
.I1(p_s2_o13_2),
.I2(p_s2_o13_3),
.I3(p_s2_o13_4),
.I4(p_s2_o13_5),
.I5(p_s2_o14_0));

wire p_s3_o15_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o13_t86_z2_v0 (
.O6(p_s3_o15_0),
.O5(),
.I0(p_s2_o13_1),
.I1(p_s2_o13_2),
.I2(p_s2_o13_3),
.I3(p_s2_o13_4),
.I4(p_s2_o13_5),
.I5(p_s2_o14_0));

/////////STEP3----ORDER14////////////

wire p_s3_o15_1;
wire p_s3_o14_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o14_t67_z0_v0 (
.O6(p_s3_o15_1),
.O5(p_s3_o14_2),
.I0(p_s2_o14_1),
.I1(p_s2_o14_2),
.I2(p_s2_o14_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER15////////////

wire p_s3_o15_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o15_t87_z0_v0 (
.O6(p_s3_o15_2),
.O5(),
.I0(p_s2_o15_0),
.I1(p_s2_o15_1),
.I2(p_s2_o15_2),
.I3(p_s2_o15_3),
.I4(p_s2_o15_4),
.I5(p_s2_o16_0));

wire p_s3_o16_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o15_t87_z1_v0 (
.O6(p_s3_o16_0),
.O5(),
.I0(p_s2_o15_0),
.I1(p_s2_o15_1),
.I2(p_s2_o15_2),
.I3(p_s2_o15_3),
.I4(p_s2_o15_4),
.I5(p_s2_o16_0));

wire p_s3_o17_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o15_t87_z2_v0 (
.O6(p_s3_o17_0),
.O5(),
.I0(p_s2_o15_0),
.I1(p_s2_o15_1),
.I2(p_s2_o15_2),
.I3(p_s2_o15_3),
.I4(p_s2_o15_4),
.I5(p_s2_o16_0));

/////////STEP3----ORDER16////////////

wire p_s3_o16_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o16_t88_z0_v0 (
.O6(p_s3_o16_1),
.O5(),
.I0(p_s2_o16_1),
.I1(p_s2_o16_2),
.I2(p_s2_o16_3),
.I3(p_s2_o16_4),
.I4(p_s2_o16_5),
.I5(p_s2_o17_0));

wire p_s3_o17_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o16_t88_z1_v0 (
.O6(p_s3_o17_1),
.O5(),
.I0(p_s2_o16_1),
.I1(p_s2_o16_2),
.I2(p_s2_o16_3),
.I3(p_s2_o16_4),
.I4(p_s2_o16_5),
.I5(p_s2_o17_0));

wire p_s3_o18_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o16_t88_z2_v0 (
.O6(p_s3_o18_0),
.O5(),
.I0(p_s2_o16_1),
.I1(p_s2_o16_2),
.I2(p_s2_o16_3),
.I3(p_s2_o16_4),
.I4(p_s2_o16_5),
.I5(p_s2_o17_0));

/////////STEP3----ORDER17////////////

wire p_s3_o17_2;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o17_t89_z0_v0 (
.O6(p_s3_o17_2),
.O5(),
.I0(p_s2_o17_1),
.I1(p_s2_o17_2),
.I2(p_s2_o17_3),
.I3(p_s2_o17_4),
.I4(p_s2_o17_5),
.I5(p_s2_o18_0));

wire p_s3_o18_1;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o17_t89_z1_v0 (
.O6(p_s3_o18_1),
.O5(),
.I0(p_s2_o17_1),
.I1(p_s2_o17_2),
.I2(p_s2_o17_3),
.I3(p_s2_o17_4),
.I4(p_s2_o17_5),
.I5(p_s2_o18_0));

wire p_s3_o19_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o17_t89_z2_v0 (
.O6(p_s3_o19_0),
.O5(),
.I0(p_s2_o17_1),
.I1(p_s2_o17_2),
.I2(p_s2_o17_3),
.I3(p_s2_o17_4),
.I4(p_s2_o17_5),
.I5(p_s2_o18_0));

/////////STEP3----ORDER18////////////

wire p_s3_o19_1;
wire p_s3_o18_2;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o18_t68_z0_v0 (
.O6(p_s3_o19_1),
.O5(p_s3_o18_2),
.I0(p_s2_o18_1),
.I1(p_s2_o18_2),
.I2(p_s2_o18_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o19_2;
wire p_s3_o18_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o18_t77_z0_v0 (
.O6(p_s3_o19_2),
.O5(p_s3_o18_3),
.I0(a[7]),
.I1(b[14]),
.I2(a[6]),
.I3(b[15]),
.I4(p_s2_o18_4),
.I5(1'b1));

/////////STEP3----ORDER19////////////

wire p_s3_o19_3;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s3_o19_t90_z0_v0 (
.O6(p_s3_o19_3),
.O5(),
.I0(p_s2_o19_0),
.I1(p_s2_o19_1),
.I2(p_s2_o19_2),
.I3(p_s1_o19_1),
.I4(p_s1_o19_2),
.I5(p_s2_o20_0));

wire p_s3_o20_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s3_o19_t90_z1_v0 (
.O6(p_s3_o20_0),
.O5(),
.I0(p_s2_o19_0),
.I1(p_s2_o19_1),
.I2(p_s2_o19_2),
.I3(p_s1_o19_1),
.I4(p_s1_o19_2),
.I5(p_s2_o20_0));

wire p_s3_o21_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s3_o19_t90_z2_v0 (
.O6(p_s3_o21_0),
.O5(),
.I0(p_s2_o19_0),
.I1(p_s2_o19_1),
.I2(p_s2_o19_2),
.I3(p_s1_o19_1),
.I4(p_s1_o19_2),
.I5(p_s2_o20_0));

/////////STEP3----ORDER20////////////

wire p_s3_o21_1;
wire p_s3_o20_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s3_o20_t69_z0_v0 (
.O6(p_s3_o21_1),
.O5(p_s3_o20_1),
.I0(p_s2_o20_1),
.I1(p_s2_o20_2),
.I2(p_s2_o20_3),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER21////////////

wire p_s3_o22_0;
wire p_s3_o21_2;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o21_t71_z0_v0 (
.O6(p_s3_o22_0),
.O5(p_s3_o21_2),
.I0(a[13]),
.I1(b[11]),
.I2(p_s2_o21_0),
.I3(p_s2_o21_1),
.I4(1'b0),
.I5(1'b1));

wire p_s3_o22_1;
wire p_s3_o21_3;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o21_t78_z0_v0 (
.O6(p_s3_o22_1),
.O5(p_s3_o21_3),
.I0(a[12]),
.I1(b[12]),
.I2(a[11]),
.I3(b[13]),
.I4(p_s2_o21_2),
.I5(1'b1));

wire p_s3_o22_2;
wire p_s3_o21_4;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o21_t78_z0_v1 (
.O6(p_s3_o22_2),
.O5(p_s3_o21_4),
.I0(a[10]),
.I1(b[14]),
.I2(a[9]),
.I3(b[15]),
.I4(p_s2_o21_3),
.I5(1'b1));

/////////STEP3----ORDER22////////////

wire p_s3_o23_0;
wire p_s3_o22_3;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o22_t72_z0_v0 (
.O6(p_s3_o23_0),
.O5(p_s3_o22_3),
.I0(a[10]),
.I1(b[15]),
.I2(p_s2_o22_0),
.I3(p_s1_o22_0),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER23////////////

wire p_s3_o24_0;
wire p_s3_o23_1;
LUT6_2 #(
.INIT(64'hF880F88087788778)
) LUT6_2_inst_s3_o23_t73_z0_v0 (
.O6(p_s3_o24_0),
.O5(p_s3_o23_1),
.I0(a[11]),
.I1(b[15]),
.I2(p_s2_o23_0),
.I3(p_s1_o23_1),
.I4(1'b0),
.I5(1'b1));

/////////STEP3----ORDER24////////////

wire p_s3_o25_0;
wire p_s3_o24_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o24_t79_z0_v0 (
.O6(p_s3_o25_0),
.O5(p_s3_o24_1),
.I0(a[13]),
.I1(b[14]),
.I2(a[12]),
.I3(b[15]),
.I4(p_s2_o24_0),
.I5(1'b1));

/////////STEP3----ORDER25////////////

wire p_s3_o26_0;
wire p_s3_o25_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s3_o25_t80_z0_v0 (
.O6(p_s3_o26_0),
.O5(p_s3_o25_1),
.I0(a[15]),
.I1(b[13]),
.I2(a[14]),
.I3(b[14]),
.I4(p_s2_o25_0),
.I5(1'b1));

/////////STEP3----ORDER26////////////

/////////STEP3----ORDER27////////////

/////////STEP4----ORDER0////////////

LUT6_2 #(
.INIT(64'h8778877808800880)
) LUT6_2_inst_oo0 (
.O6(P[0]),
.O5(G[0]),
.I0(a[0]),
.I1(b[3]),
.I2(C0),
.I3(p_s0_o0_0),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER1////////////

LUT6_2 #(
.INIT(64'h8778787878000000)
) LUT6_2_inst_oo1 (
.O6(P[1]),
.O5(G[1]),
.I0(a[0]),
.I1(b[4]),
.I2(p_s2_o1_0),
.I3(C0),
.I4(p_s0_o0_0),
.I5(1'b1));

/////////STEP4----ORDER2////////////

LUT6_2 #(
.INIT(64'h9666666660000000)
) LUT6_2_inst_oo2 (
.O6(P[2]),
.O5(G[2]),
.I0(p_s3_o2_0),
.I1(p_s3_o2_1),
.I2(a[0]),
.I3(b[4]),
.I4(p_s2_o1_0),
.I5(1'b1));

/////////STEP4----ORDER3////////////

wire p_s4_o4_0;
wire p_s4_o3_0;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o3_t101_z0_v0 (
.O6(p_s4_o4_0),
.O5(p_s4_o3_0),
.I0(p_s3_o3_0),
.I1(p_s3_o3_1),
.I2(p_s2_o3_0),
.I3(p_s3_o4_0),
.I4(p_s2_o4_1),
.I5(1'b1));

wire p_s4_o5_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o3_t101_z1_v0 (
.O6(p_s4_o5_0),
.O5(),
.I0(p_s3_o3_0),
.I1(p_s3_o3_1),
.I2(p_s2_o3_0),
.I3(p_s3_o4_0),
.I4(p_s2_o4_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo3 (
.O6(P[3]),
.O5(G[3]),
.I0(p_s4_o3_0),
.I1(p_s2_o3_1),
.I2(p_s3_o2_0),
.I3(p_s3_o2_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER4////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo4 (
.O6(P[4]),
.O5(G[4]),
.I0(p_s4_o4_0),
.I1(p_s2_o4_2),
.I2(p_s4_o3_0),
.I3(p_s2_o3_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER5////////////

wire p_s4_o5_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o5_t96_z0_v0 (
.O6(p_s4_o5_1),
.O5(),
.I0(p_s3_o5_0),
.I1(p_s2_o5_0),
.I2(p_s2_o5_1),
.I3(p_s2_o5_2),
.I4(p_s2_o5_3),
.I5(p_s3_o6_0));

wire p_s4_o6_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o5_t96_z1_v0 (
.O6(p_s4_o6_0),
.O5(),
.I0(p_s3_o5_0),
.I1(p_s2_o5_0),
.I2(p_s2_o5_1),
.I3(p_s2_o5_2),
.I4(p_s2_o5_3),
.I5(p_s3_o6_0));

wire p_s4_o7_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o5_t96_z2_v0 (
.O6(p_s4_o7_0),
.O5(),
.I0(p_s3_o5_0),
.I1(p_s2_o5_0),
.I2(p_s2_o5_1),
.I3(p_s2_o5_2),
.I4(p_s2_o5_3),
.I5(p_s3_o6_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo5 (
.O6(P[5]),
.O5(G[5]),
.I0(p_s4_o5_0),
.I1(p_s4_o5_1),
.I2(p_s4_o4_0),
.I3(p_s2_o4_2),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER6////////////

LUT6_2 #(
.INIT(64'h8778787878000000)
) LUT6_2_inst_oo6 (
.O6(P[6]),
.O5(G[6]),
.I0(a[0]),
.I1(b[9]),
.I2(p_s4_o6_0),
.I3(p_s4_o5_0),
.I4(p_s4_o5_1),
.I5(1'b1));

/////////STEP4----ORDER7////////////

wire p_s4_o8_0;
wire p_s4_o7_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s4_o7_t91_z0_v0 (
.O6(p_s4_o8_0),
.O5(p_s4_o7_1),
.I0(p_s3_o7_0),
.I1(p_s3_o7_1),
.I2(p_s3_o7_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666666660000000)
) LUT6_2_inst_oo7 (
.O6(P[7]),
.O5(G[7]),
.I0(p_s4_o7_0),
.I1(p_s4_o7_1),
.I2(a[0]),
.I3(b[9]),
.I4(p_s4_o6_0),
.I5(1'b1));

/////////STEP4----ORDER8////////////

wire p_s4_o8_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o8_t97_z0_v0 (
.O6(p_s4_o8_1),
.O5(),
.I0(p_s3_o8_0),
.I1(p_s3_o8_1),
.I2(p_s3_o8_2),
.I3(p_s3_o8_3),
.I4(p_s0_o8_1),
.I5(p_s3_o9_0));

wire p_s4_o9_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o8_t97_z1_v0 (
.O6(p_s4_o9_0),
.O5(),
.I0(p_s3_o8_0),
.I1(p_s3_o8_1),
.I2(p_s3_o8_2),
.I3(p_s3_o8_3),
.I4(p_s0_o8_1),
.I5(p_s3_o9_0));

wire p_s4_o10_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o8_t97_z2_v0 (
.O6(p_s4_o10_0),
.O5(),
.I0(p_s3_o8_0),
.I1(p_s3_o8_1),
.I2(p_s3_o8_2),
.I3(p_s3_o8_3),
.I4(p_s0_o8_1),
.I5(p_s3_o9_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo8 (
.O6(P[8]),
.O5(G[8]),
.I0(p_s4_o8_0),
.I1(p_s4_o8_1),
.I2(p_s4_o7_0),
.I3(p_s4_o7_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER9////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo9 (
.O6(P[9]),
.O5(G[9]),
.I0(p_s4_o9_0),
.I1(p_s3_o9_1),
.I2(p_s4_o8_0),
.I3(p_s4_o8_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER10////////////

wire p_s4_o11_0;
wire p_s4_o10_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s4_o10_t92_z0_v0 (
.O6(p_s4_o11_0),
.O5(p_s4_o10_1),
.I0(p_s3_o10_0),
.I1(p_s3_o10_1),
.I2(p_s3_o10_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo10 (
.O6(P[10]),
.O5(G[10]),
.I0(p_s4_o10_0),
.I1(p_s4_o10_1),
.I2(p_s4_o9_0),
.I3(p_s3_o9_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER11////////////

wire p_s4_o11_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o11_t98_z0_v0 (
.O6(p_s4_o11_1),
.O5(),
.I0(p_s3_o11_0),
.I1(p_s3_o11_1),
.I2(p_s3_o11_2),
.I3(p_s3_o11_3),
.I4(p_s2_o11_7),
.I5(p_s3_o12_0));

wire p_s4_o12_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o11_t98_z1_v0 (
.O6(p_s4_o12_0),
.O5(),
.I0(p_s3_o11_0),
.I1(p_s3_o11_1),
.I2(p_s3_o11_2),
.I3(p_s3_o11_3),
.I4(p_s2_o11_7),
.I5(p_s3_o12_0));

wire p_s4_o13_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o11_t98_z2_v0 (
.O6(p_s4_o13_0),
.O5(),
.I0(p_s3_o11_0),
.I1(p_s3_o11_1),
.I2(p_s3_o11_2),
.I3(p_s3_o11_3),
.I4(p_s2_o11_7),
.I5(p_s3_o12_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo11 (
.O6(P[11]),
.O5(G[11]),
.I0(p_s4_o11_0),
.I1(p_s4_o11_1),
.I2(p_s4_o10_0),
.I3(p_s4_o10_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER12////////////

wire p_s4_o13_1;
wire p_s4_o12_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o12_t102_z0_v0 (
.O6(p_s4_o13_1),
.O5(p_s4_o12_1),
.I0(p_s3_o12_1),
.I1(p_s3_o12_2),
.I2(p_s3_o12_3),
.I3(p_s3_o13_0),
.I4(p_s3_o13_1),
.I5(1'b1));

wire p_s4_o14_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o12_t102_z1_v0 (
.O6(p_s4_o14_0),
.O5(),
.I0(p_s3_o12_1),
.I1(p_s3_o12_2),
.I2(p_s3_o12_3),
.I3(p_s3_o13_0),
.I4(p_s3_o13_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo12 (
.O6(P[12]),
.O5(G[12]),
.I0(p_s4_o12_0),
.I1(p_s4_o12_1),
.I2(p_s4_o11_0),
.I3(p_s4_o11_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER13////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo13 (
.O6(P[13]),
.O5(G[13]),
.I0(p_s4_o13_0),
.I1(p_s4_o13_1),
.I2(p_s4_o12_0),
.I3(p_s4_o12_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER14////////////

wire p_s4_o14_1;
LUT6_2 #(
.INIT(64'h6996966996696996)
) LUT6_2_inst_s4_o14_t95_z0_v0 (
.O6(p_s4_o14_1),
.O5(),
.I0(p_s3_o14_0),
.I1(p_s3_o14_1),
.I2(p_s3_o14_2),
.I3(p_s2_o14_4),
.I4(p_s2_o14_5),
.I5(p_s2_o14_6));

wire p_s4_o15_0;
LUT6_2 #(
.INIT(64'h8117177E177E7EE8)
) LUT6_2_inst_s4_o14_t95_z1_v0 (
.O6(p_s4_o15_0),
.O5(),
.I0(p_s3_o14_0),
.I1(p_s3_o14_1),
.I2(p_s3_o14_2),
.I3(p_s2_o14_4),
.I4(p_s2_o14_5),
.I5(p_s2_o14_6));

wire p_s4_o16_0;
LUT6_2 #(
.INIT(64'hFEE8E880E8808000)
) LUT6_2_inst_s4_o14_t95_z2_v0 (
.O6(p_s4_o16_0),
.O5(),
.I0(p_s3_o14_0),
.I1(p_s3_o14_1),
.I2(p_s3_o14_2),
.I3(p_s2_o14_4),
.I4(p_s2_o14_5),
.I5(p_s2_o14_6));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo14 (
.O6(P[14]),
.O5(G[14]),
.I0(p_s4_o14_0),
.I1(p_s4_o14_1),
.I2(p_s4_o13_0),
.I3(p_s4_o13_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER15////////////

wire p_s4_o16_1;
wire p_s4_o15_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o15_t103_z0_v0 (
.O6(p_s4_o16_1),
.O5(p_s4_o15_1),
.I0(p_s3_o15_0),
.I1(p_s3_o15_1),
.I2(p_s3_o15_2),
.I3(p_s3_o16_0),
.I4(p_s3_o16_1),
.I5(1'b1));

wire p_s4_o17_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o15_t103_z1_v0 (
.O6(p_s4_o17_0),
.O5(),
.I0(p_s3_o15_0),
.I1(p_s3_o15_1),
.I2(p_s3_o15_2),
.I3(p_s3_o16_0),
.I4(p_s3_o16_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo15 (
.O6(P[15]),
.O5(G[15]),
.I0(p_s4_o15_0),
.I1(p_s4_o15_1),
.I2(p_s4_o14_0),
.I3(p_s4_o14_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER16////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo16 (
.O6(P[16]),
.O5(G[16]),
.I0(p_s4_o16_0),
.I1(p_s4_o16_1),
.I2(p_s4_o15_0),
.I3(p_s4_o15_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER17////////////

wire p_s4_o18_0;
wire p_s4_o17_1;
LUT6_2 #(
.INIT(64'hE8E8E8E896969696)
) LUT6_2_inst_s4_o17_t93_z0_v0 (
.O6(p_s4_o18_0),
.O5(p_s4_o17_1),
.I0(p_s3_o17_0),
.I1(p_s3_o17_1),
.I2(p_s3_o17_2),
.I3(1'b0),
.I4(1'b0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo17 (
.O6(P[17]),
.O5(G[17]),
.I0(p_s4_o17_0),
.I1(p_s4_o17_1),
.I2(p_s4_o16_0),
.I3(p_s4_o16_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER18////////////

wire p_s4_o18_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o18_t99_z0_v0 (
.O6(p_s4_o18_1),
.O5(),
.I0(p_s3_o18_0),
.I1(p_s3_o18_1),
.I2(p_s3_o18_2),
.I3(p_s3_o18_3),
.I4(p_s2_o18_5),
.I5(p_s3_o19_0));

wire p_s4_o19_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o18_t99_z1_v0 (
.O6(p_s4_o19_0),
.O5(),
.I0(p_s3_o18_0),
.I1(p_s3_o18_1),
.I2(p_s3_o18_2),
.I3(p_s3_o18_3),
.I4(p_s2_o18_5),
.I5(p_s3_o19_0));

wire p_s4_o20_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o18_t99_z2_v0 (
.O6(p_s4_o20_0),
.O5(),
.I0(p_s3_o18_0),
.I1(p_s3_o18_1),
.I2(p_s3_o18_2),
.I3(p_s3_o18_3),
.I4(p_s2_o18_5),
.I5(p_s3_o19_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo18 (
.O6(P[18]),
.O5(G[18]),
.I0(p_s4_o18_0),
.I1(p_s4_o18_1),
.I2(p_s4_o17_0),
.I3(p_s4_o17_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER19////////////

wire p_s4_o20_1;
wire p_s4_o19_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o19_t104_z0_v0 (
.O6(p_s4_o20_1),
.O5(p_s4_o19_1),
.I0(p_s3_o19_1),
.I1(p_s3_o19_2),
.I2(p_s3_o19_3),
.I3(p_s3_o20_0),
.I4(p_s3_o20_1),
.I5(1'b1));

wire p_s4_o21_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o19_t104_z1_v0 (
.O6(p_s4_o21_0),
.O5(),
.I0(p_s3_o19_1),
.I1(p_s3_o19_2),
.I2(p_s3_o19_3),
.I3(p_s3_o20_0),
.I4(p_s3_o20_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo19 (
.O6(P[19]),
.O5(G[19]),
.I0(p_s4_o19_0),
.I1(p_s4_o19_1),
.I2(p_s4_o18_0),
.I3(p_s4_o18_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER20////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo20 (
.O6(P[20]),
.O5(G[20]),
.I0(p_s4_o20_0),
.I1(p_s4_o20_1),
.I2(p_s4_o19_0),
.I3(p_s4_o19_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER21////////////

wire p_s4_o21_1;
LUT6_2 #(
.INIT(64'h9669699696696996)
) LUT6_2_inst_s4_o21_t100_z0_v0 (
.O6(p_s4_o21_1),
.O5(),
.I0(p_s3_o21_0),
.I1(p_s3_o21_1),
.I2(p_s3_o21_2),
.I3(p_s3_o21_3),
.I4(p_s3_o21_4),
.I5(p_s3_o22_0));

wire p_s4_o22_0;
LUT6_2 #(
.INIT(64'hE8818117177E7EE8)
) LUT6_2_inst_s4_o21_t100_z1_v0 (
.O6(p_s4_o22_0),
.O5(),
.I0(p_s3_o21_0),
.I1(p_s3_o21_1),
.I2(p_s3_o21_2),
.I3(p_s3_o21_3),
.I4(p_s3_o21_4),
.I5(p_s3_o22_0));

wire p_s4_o23_0;
LUT6_2 #(
.INIT(64'hFFFEFEE8E8808000)
) LUT6_2_inst_s4_o21_t100_z2_v0 (
.O6(p_s4_o23_0),
.O5(),
.I0(p_s3_o21_0),
.I1(p_s3_o21_1),
.I2(p_s3_o21_2),
.I3(p_s3_o21_3),
.I4(p_s3_o21_4),
.I5(p_s3_o22_0));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo21 (
.O6(P[21]),
.O5(G[21]),
.I0(p_s4_o21_0),
.I1(p_s4_o21_1),
.I2(p_s4_o20_0),
.I3(p_s4_o20_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER22////////////

wire p_s4_o23_1;
wire p_s4_o22_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o22_t105_z0_v0 (
.O6(p_s4_o23_1),
.O5(p_s4_o22_1),
.I0(p_s3_o22_1),
.I1(p_s3_o22_2),
.I2(p_s3_o22_3),
.I3(p_s3_o23_0),
.I4(p_s3_o23_1),
.I5(1'b1));

wire p_s4_o24_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o22_t105_z1_v0 (
.O6(p_s4_o24_0),
.O5(),
.I0(p_s3_o22_1),
.I1(p_s3_o22_2),
.I2(p_s3_o22_3),
.I3(p_s3_o23_0),
.I4(p_s3_o23_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo22 (
.O6(P[22]),
.O5(G[22]),
.I0(p_s4_o22_0),
.I1(p_s4_o22_1),
.I2(p_s4_o21_0),
.I3(p_s4_o21_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER23////////////

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo23 (
.O6(P[23]),
.O5(G[23]),
.I0(p_s4_o23_0),
.I1(p_s4_o23_1),
.I2(p_s4_o22_0),
.I3(p_s4_o22_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER24////////////

wire p_s4_o25_0;
wire p_s4_o24_1;
LUT6_2 #(
.INIT(64'hE81717E896969696)
) LUT6_2_inst_s4_o24_t106_z0_v0 (
.O6(p_s4_o25_0),
.O5(p_s4_o24_1),
.I0(p_s3_o24_0),
.I1(p_s3_o24_1),
.I2(p_s2_o24_1),
.I3(p_s3_o25_0),
.I4(p_s3_o25_1),
.I5(1'b1));

wire p_s4_o26_0;
LUT6_2 #(
.INIT(64'hFFE8E800FFE8E800)
) LUT6_2_inst_s4_o24_t106_z1_v0 (
.O6(p_s4_o26_0),
.O5(),
.I0(p_s3_o24_0),
.I1(p_s3_o24_1),
.I2(p_s2_o24_1),
.I3(p_s3_o25_0),
.I4(p_s3_o25_1),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666966660006000)
) LUT6_2_inst_oo24 (
.O6(P[24]),
.O5(G[24]),
.I0(p_s4_o24_0),
.I1(p_s4_o24_1),
.I2(p_s4_o23_0),
.I3(p_s4_o23_1),
.I4(1'b1),
.I5(1'b1));

/////////STEP4----ORDER25////////////

LUT6_2 #(
.INIT(64'h8778787878000000)
) LUT6_2_inst_oo25 (
.O6(P[25]),
.O5(G[25]),
.I0(a[13]),
.I1(b[15]),
.I2(p_s4_o25_0),
.I3(p_s4_o24_0),
.I4(p_s4_o24_1),
.I5(1'b1));

/////////STEP4----ORDER26////////////

wire p_s4_o27_0;
wire p_s4_o26_1;
LUT6_2 #(
.INIT(64'hF888800087777888)
) LUT6_2_inst_s4_o26_t94_z0_v0 (
.O6(p_s4_o27_0),
.O5(p_s4_o26_1),
.I0(a[15]),
.I1(b[14]),
.I2(a[14]),
.I3(b[15]),
.I4(p_s3_o26_0),
.I5(1'b1));

LUT6_2 #(
.INIT(64'h9666666660000000)
) LUT6_2_inst_oo26 (
.O6(P[26]),
.O5(G[26]),
.I0(p_s4_o26_0),
.I1(p_s4_o26_1),
.I2(a[13]),
.I3(b[15]),
.I4(p_s4_o25_0),
.I5(1'b1));

/////////STEP4----ORDER27////////////

LUT6_2 #(
.INIT(64'h87777888F8888000)
) LUT6_2_inst_ooo (
.O6(P[27]),
.O5(G[27]),
.I0(b[15]),
.I1(a[15]),
.I2(p_s4_o26_0),
.I3(p_s4_o26_1),
.I4(p_s4_o27_0),
.I5(1'b1));

wire [3:0] carry_o_0;
CARRY4  CARRY4_inst_0(
.CO(carry_o_0),
.O(r[6:3]),
.CI(C1),
.CYINIT(1'b0),
.DI(G[3:0]),
.S(P[3:0]));

wire [3:0] carry_o_1;
CARRY4  CARRY4_inst_1(
.CO(carry_o_1),
.O(r[10:7]),
.CI(carry_o_0[3]),
.CYINIT(1'b0),
.DI(G[7:4]),
.S(P[7:4]));

wire [3:0] carry_o_2;
CARRY4  CARRY4_inst_2(
.CO(carry_o_2),
.O(r[14:11]),
.CI(carry_o_1[3]),
.CYINIT(1'b0),
.DI(G[11:8]),
.S(P[11:8]));

wire [3:0] carry_o_3;
CARRY4  CARRY4_inst_3(
.CO(carry_o_3),
.O(r[18:15]),
.CI(carry_o_2[3]),
.CYINIT(1'b0),
.DI(G[15:12]),
.S(P[15:12]));

wire [3:0] carry_o_4;
CARRY4  CARRY4_inst_4(
.CO(carry_o_4),
.O(r[22:19]),
.CI(carry_o_3[3]),
.CYINIT(1'b0),
.DI(G[19:16]),
.S(P[19:16]));

wire [3:0] carry_o_5;
CARRY4  CARRY4_inst_5(
.CO(carry_o_5),
.O(r[26:23]),
.CI(carry_o_4[3]),
.CYINIT(1'b0),
.DI(G[23:20]),
.S(P[23:20]));

wire [3:0] carry_o_6;
CARRY4  CARRY4_inst_6(
.CO(carry_o_6),
.O(r[30:27]),
.CI(carry_o_5[3]),
.CYINIT(1'b0),
.DI(G[27:24]),
.S(P[27:24]));

assign  r[31] = carry_o_6[3] | (P[27] & G[27]);
//v2024-09-29 04:44:44.798719
endmodule
